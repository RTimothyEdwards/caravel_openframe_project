magic
tech sky130A
magscale 1 2
timestamp 1685879372
<< viali >>
rect 4261 13413 4295 13447
rect 4721 13413 4755 13447
rect 8493 13413 8527 13447
rect 9045 13413 9079 13447
rect 13093 13413 13127 13447
rect 13369 13413 13403 13447
rect 16359 13413 16393 13447
rect 3893 13345 3927 13379
rect 6561 13345 6595 13379
rect 9643 13345 9677 13379
rect 17325 13345 17359 13379
rect 4905 13277 4939 13311
rect 5549 13277 5583 13311
rect 5703 13277 5737 13311
rect 6745 13277 6779 13311
rect 7021 13277 7055 13311
rect 8125 13277 8159 13311
rect 9229 13277 9263 13311
rect 9540 13277 9574 13311
rect 10241 13277 10275 13311
rect 10333 13277 10367 13311
rect 12056 13277 12090 13311
rect 12725 13277 12759 13311
rect 13553 13277 13587 13311
rect 14197 13277 14231 13311
rect 15577 13277 15611 13311
rect 16288 13277 16322 13311
rect 16773 13277 16807 13311
rect 17785 13277 17819 13311
rect 5917 13209 5951 13243
rect 7389 13209 7423 13243
rect 14657 13209 14691 13243
rect 14749 13209 14783 13243
rect 15761 13209 15795 13243
rect 17233 13209 17267 13243
rect 4261 13141 4295 13175
rect 6929 13141 6963 13175
rect 7481 13141 7515 13175
rect 8493 13141 8527 13175
rect 10241 13141 10275 13175
rect 12127 13141 12161 13175
rect 13093 13141 13127 13175
rect 17601 13141 17635 13175
rect 8677 12937 8711 12971
rect 13369 12937 13403 12971
rect 4353 12869 4387 12903
rect 5825 12869 5859 12903
rect 10011 12869 10045 12903
rect 10701 12869 10735 12903
rect 12081 12869 12115 12903
rect 12173 12869 12207 12903
rect 17233 12869 17267 12903
rect 3065 12801 3099 12835
rect 3617 12801 3651 12835
rect 3893 12801 3927 12835
rect 4445 12801 4479 12835
rect 6469 12801 6503 12835
rect 7021 12801 7055 12835
rect 8309 12801 8343 12835
rect 9505 12801 9539 12835
rect 9689 12801 9723 12835
rect 9781 12801 9815 12835
rect 9873 12801 9907 12835
rect 10517 12801 10551 12835
rect 10785 12801 10819 12835
rect 10931 12801 10965 12835
rect 14657 12801 14691 12835
rect 15209 12801 15243 12835
rect 15761 12801 15795 12835
rect 15945 12801 15979 12835
rect 16037 12801 16071 12835
rect 16773 12801 16807 12835
rect 17325 12801 17359 12835
rect 18036 12801 18070 12835
rect 6009 12733 6043 12767
rect 8677 12733 8711 12767
rect 10149 12733 10183 12767
rect 11621 12733 11655 12767
rect 13001 12733 13035 12767
rect 13369 12733 13403 12767
rect 15025 12733 15059 12767
rect 3617 12665 3651 12699
rect 7021 12665 7055 12699
rect 15577 12665 15611 12699
rect 11069 12597 11103 12631
rect 18107 12597 18141 12631
rect 9965 12393 9999 12427
rect 13185 12393 13219 12427
rect 13737 12393 13771 12427
rect 15163 12393 15197 12427
rect 16037 12393 16071 12427
rect 17693 12393 17727 12427
rect 2697 12325 2731 12359
rect 4629 12325 4663 12359
rect 7757 12325 7791 12359
rect 3065 12257 3099 12291
rect 4169 12257 4203 12291
rect 7297 12257 7331 12291
rect 7849 12257 7883 12291
rect 8217 12257 8251 12291
rect 11069 12257 11103 12291
rect 17693 12257 17727 12291
rect 1869 12189 1903 12223
rect 2145 12189 2179 12223
rect 3249 12189 3283 12223
rect 3525 12189 3559 12223
rect 5032 12189 5066 12223
rect 6285 12189 6319 12223
rect 6653 12189 6687 12223
rect 8401 12189 8435 12223
rect 8677 12189 8711 12223
rect 9229 12189 9263 12223
rect 9413 12189 9447 12223
rect 10241 12189 10275 12223
rect 10701 12189 10735 12223
rect 11253 12189 11287 12223
rect 12173 12189 12207 12223
rect 12633 12189 12667 12223
rect 13001 12189 13035 12223
rect 13645 12189 13679 12223
rect 14197 12189 14231 12223
rect 14565 12189 14599 12223
rect 15060 12189 15094 12223
rect 15485 12189 15519 12223
rect 16037 12189 16071 12223
rect 17325 12189 17359 12223
rect 18245 12189 18279 12223
rect 2513 12121 2547 12155
rect 4721 12121 4755 12155
rect 5135 12121 5169 12155
rect 9965 12121 9999 12155
rect 12817 12121 12851 12155
rect 12909 12121 12943 12155
rect 1685 12053 1719 12087
rect 2053 12053 2087 12087
rect 3433 12053 3467 12087
rect 6653 12053 6687 12087
rect 8585 12053 8619 12087
rect 9321 12053 9355 12087
rect 10149 12053 10183 12087
rect 12357 12053 12391 12087
rect 14565 12053 14599 12087
rect 18337 12053 18371 12087
rect 4629 11849 4663 11883
rect 5917 11849 5951 11883
rect 8033 11849 8067 11883
rect 12817 11849 12851 11883
rect 14013 11849 14047 11883
rect 14841 11849 14875 11883
rect 8493 11781 8527 11815
rect 12449 11781 12483 11815
rect 1501 11713 1535 11747
rect 2053 11713 2087 11747
rect 3525 11713 3559 11747
rect 4445 11713 4479 11747
rect 4721 11713 4755 11747
rect 5089 11713 5123 11747
rect 6101 11713 6135 11747
rect 7389 11713 7423 11747
rect 7849 11713 7883 11747
rect 8125 11713 8159 11747
rect 8677 11713 8711 11747
rect 8861 11713 8895 11747
rect 9873 11713 9907 11747
rect 9965 11713 9999 11747
rect 10057 11713 10091 11747
rect 10241 11713 10275 11747
rect 10517 11713 10551 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 10885 11713 10919 11747
rect 11713 11713 11747 11747
rect 12265 11713 12299 11747
rect 12541 11713 12575 11747
rect 12633 11713 12667 11747
rect 13093 11713 13127 11747
rect 13645 11713 13679 11747
rect 15025 11713 15059 11747
rect 16405 11713 16439 11747
rect 16865 11713 16899 11747
rect 17417 11713 17451 11747
rect 5273 11645 5307 11679
rect 7021 11645 7055 11679
rect 8953 11645 8987 11679
rect 14013 11645 14047 11679
rect 7205 11577 7239 11611
rect 7665 11577 7699 11611
rect 11069 11577 11103 11611
rect 2053 11509 2087 11543
rect 3341 11509 3375 11543
rect 4261 11509 4295 11543
rect 9597 11509 9631 11543
rect 11805 11509 11839 11543
rect 13185 11509 13219 11543
rect 16221 11509 16255 11543
rect 17417 11509 17451 11543
rect 4629 11305 4663 11339
rect 6653 11305 6687 11339
rect 8125 11305 8159 11339
rect 10609 11305 10643 11339
rect 13277 11305 13311 11339
rect 9045 11237 9079 11271
rect 10149 11237 10183 11271
rect 18153 11237 18187 11271
rect 1777 11169 1811 11203
rect 7021 11169 7055 11203
rect 8585 11169 8619 11203
rect 8677 11169 8711 11203
rect 9505 11169 9539 11203
rect 11529 11169 11563 11203
rect 12633 11169 12667 11203
rect 14565 11169 14599 11203
rect 15577 11169 15611 11203
rect 17785 11169 17819 11203
rect 2973 11101 3007 11135
rect 3525 11101 3559 11135
rect 4077 11101 4111 11135
rect 4629 11101 4663 11135
rect 5984 11101 6018 11135
rect 6837 11101 6871 11135
rect 7113 11101 7147 11135
rect 8125 11101 8159 11135
rect 8381 11101 8415 11135
rect 9045 11101 9079 11135
rect 9229 11101 9263 11135
rect 9781 11101 9815 11135
rect 9965 11101 9999 11135
rect 10241 11101 10275 11135
rect 10885 11101 10919 11135
rect 10977 11101 11011 11135
rect 11069 11101 11103 11135
rect 11253 11101 11287 11135
rect 11713 11101 11747 11135
rect 11897 11101 11931 11135
rect 12265 11101 12299 11135
rect 12358 11101 12392 11135
rect 14749 11101 14783 11135
rect 14933 11101 14967 11135
rect 15209 11101 15243 11135
rect 15761 11101 15795 11135
rect 16037 11101 16071 11135
rect 16405 11101 16439 11135
rect 16957 11101 16991 11135
rect 2237 11033 2271 11067
rect 2329 11033 2363 11067
rect 3433 11033 3467 11067
rect 9873 11033 9907 11067
rect 13093 11033 13127 11067
rect 14841 11033 14875 11067
rect 15071 11033 15105 11067
rect 16865 11033 16899 11067
rect 6055 10965 6089 10999
rect 8493 10965 8527 10999
rect 13293 10965 13327 10999
rect 13461 10965 13495 10999
rect 15945 10965 15979 10999
rect 18153 10965 18187 10999
rect 2375 10761 2409 10795
rect 3249 10761 3283 10795
rect 8677 10761 8711 10795
rect 10149 10761 10183 10795
rect 10425 10761 10459 10795
rect 11897 10761 11931 10795
rect 12817 10761 12851 10795
rect 13921 10761 13955 10795
rect 16221 10761 16255 10795
rect 17233 10761 17267 10795
rect 4997 10693 5031 10727
rect 6745 10693 6779 10727
rect 15117 10693 15151 10727
rect 15210 10693 15244 10727
rect 15347 10693 15381 10727
rect 15853 10693 15887 10727
rect 18153 10693 18187 10727
rect 18245 10693 18279 10727
rect 16083 10659 16117 10693
rect 2304 10625 2338 10659
rect 3249 10625 3283 10659
rect 4445 10625 4479 10659
rect 4905 10625 4939 10659
rect 5340 10625 5374 10659
rect 6561 10625 6595 10659
rect 6837 10625 6871 10659
rect 6929 10625 6963 10659
rect 7633 10625 7667 10659
rect 7757 10625 7791 10659
rect 8953 10625 8987 10659
rect 9045 10625 9079 10659
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 10610 10625 10644 10659
rect 10701 10625 10735 10659
rect 10977 10625 11011 10659
rect 12081 10625 12115 10659
rect 12265 10625 12299 10659
rect 12357 10625 12391 10659
rect 12725 10625 12759 10659
rect 13185 10625 13219 10659
rect 13369 10625 13403 10659
rect 13553 10625 13587 10659
rect 13737 10625 13771 10659
rect 14197 10625 14231 10659
rect 15025 10625 15059 10659
rect 17693 10625 17727 10659
rect 2881 10557 2915 10591
rect 7849 10557 7883 10591
rect 10885 10557 10919 10591
rect 13461 10557 13495 10591
rect 15485 10557 15519 10591
rect 16865 10557 16899 10591
rect 14841 10489 14875 10523
rect 17233 10489 17267 10523
rect 5411 10421 5445 10455
rect 7113 10421 7147 10455
rect 7389 10421 7423 10455
rect 14289 10421 14323 10455
rect 16037 10421 16071 10455
rect 4537 10217 4571 10251
rect 9045 10217 9079 10251
rect 9505 10217 9539 10251
rect 10149 10217 10183 10251
rect 12173 10217 12207 10251
rect 13553 10217 13587 10251
rect 15301 10217 15335 10251
rect 5273 10149 5307 10183
rect 5733 10149 5767 10183
rect 7757 10149 7791 10183
rect 7941 10149 7975 10183
rect 8401 10149 8435 10183
rect 13093 10149 13127 10183
rect 15669 10149 15703 10183
rect 17141 10149 17175 10183
rect 12817 10081 12851 10115
rect 14473 10081 14507 10115
rect 2364 10013 2398 10047
rect 4905 10013 4939 10047
rect 5917 10013 5951 10047
rect 6377 10013 6411 10047
rect 6653 10013 6687 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 9230 10013 9264 10047
rect 9381 10013 9415 10047
rect 9597 10013 9631 10047
rect 10149 10013 10183 10047
rect 10327 10013 10361 10047
rect 10609 10013 10643 10047
rect 10793 10013 10827 10047
rect 11437 10013 11471 10047
rect 11621 10013 11655 10047
rect 12081 10013 12115 10047
rect 13277 10013 13311 10047
rect 13369 10013 13403 10047
rect 13645 10013 13679 10047
rect 15209 10013 15243 10047
rect 15301 10013 15335 10047
rect 15853 10013 15887 10047
rect 16773 10013 16807 10047
rect 18061 10013 18095 10047
rect 4445 9945 4479 9979
rect 7481 9945 7515 9979
rect 12633 9945 12667 9979
rect 14289 9945 14323 9979
rect 15025 9945 15059 9979
rect 15577 9945 15611 9979
rect 15761 9945 15795 9979
rect 17141 9945 17175 9979
rect 18245 9945 18279 9979
rect 2467 9877 2501 9911
rect 5273 9877 5307 9911
rect 6193 9877 6227 9911
rect 6561 9877 6595 9911
rect 10701 9877 10735 9911
rect 11529 9877 11563 9911
rect 5917 9673 5951 9707
rect 7481 9673 7515 9707
rect 11069 9673 11103 9707
rect 12173 9673 12207 9707
rect 15393 9673 15427 9707
rect 16221 9673 16255 9707
rect 7297 9605 7331 9639
rect 8033 9605 8067 9639
rect 10701 9605 10735 9639
rect 10901 9605 10935 9639
rect 14197 9605 14231 9639
rect 14381 9605 14415 9639
rect 15853 9605 15887 9639
rect 1869 9537 1903 9571
rect 3157 9537 3191 9571
rect 3709 9537 3743 9571
rect 5549 9537 5583 9571
rect 7757 9537 7791 9571
rect 9045 9537 9079 9571
rect 9137 9537 9171 9571
rect 9321 9537 9355 9571
rect 9413 9537 9447 9571
rect 9781 9537 9815 9571
rect 11897 9537 11931 9571
rect 11989 9537 12023 9571
rect 12633 9537 12667 9571
rect 12909 9537 12943 9571
rect 13461 9537 13495 9571
rect 13553 9537 13587 9571
rect 13645 9537 13679 9571
rect 14565 9537 14599 9571
rect 14657 9537 14691 9571
rect 14841 9537 14875 9571
rect 14933 9537 14967 9571
rect 15301 9537 15335 9571
rect 16037 9537 16071 9571
rect 16313 9537 16347 9571
rect 16865 9537 16899 9571
rect 17417 9537 17451 9571
rect 2145 9469 2179 9503
rect 5917 9469 5951 9503
rect 6929 9469 6963 9503
rect 8033 9469 8067 9503
rect 10057 9469 10091 9503
rect 3709 9401 3743 9435
rect 7849 9401 7883 9435
rect 8861 9401 8895 9435
rect 12725 9401 12759 9435
rect 12817 9401 12851 9435
rect 13829 9401 13863 9435
rect 7297 9333 7331 9367
rect 9873 9333 9907 9367
rect 9965 9333 9999 9367
rect 10885 9333 10919 9367
rect 12449 9333 12483 9367
rect 17417 9333 17451 9367
rect 3065 9129 3099 9163
rect 4997 9129 5031 9163
rect 7941 9129 7975 9163
rect 9137 9129 9171 9163
rect 9781 9129 9815 9163
rect 11345 9129 11379 9163
rect 12081 9129 12115 9163
rect 16681 9129 16715 9163
rect 4353 9061 4387 9095
rect 10241 9061 10275 9095
rect 13461 9061 13495 9095
rect 14657 9061 14691 9095
rect 15485 9061 15519 9095
rect 17601 9061 17635 9095
rect 3893 8993 3927 9027
rect 4445 8993 4479 9027
rect 7297 8993 7331 9027
rect 12541 8993 12575 9027
rect 14289 8993 14323 9027
rect 15853 8993 15887 9027
rect 2053 8925 2087 8959
rect 2329 8925 2363 8959
rect 2513 8925 2547 8959
rect 3249 8925 3283 8959
rect 3525 8925 3559 8959
rect 5524 8925 5558 8959
rect 7113 8925 7147 8959
rect 7205 8925 7239 8959
rect 7401 8925 7435 8959
rect 8309 8925 8343 8959
rect 8493 8925 8527 8959
rect 9045 8925 9079 8959
rect 9689 8925 9723 8959
rect 9873 8925 9907 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 11253 8925 11287 8959
rect 11437 8925 11471 8959
rect 12449 8925 12483 8959
rect 12633 8925 12667 8959
rect 12909 8925 12943 8959
rect 13093 8925 13127 8959
rect 13369 8925 13403 8959
rect 13553 8925 13587 8959
rect 14473 8925 14507 8959
rect 14933 8925 14967 8959
rect 15117 8925 15151 8959
rect 15301 8925 15335 8959
rect 16221 8925 16255 8959
rect 16865 8925 16899 8959
rect 17141 8925 17175 8959
rect 18004 8925 18038 8959
rect 1869 8857 1903 8891
rect 4905 8857 4939 8891
rect 6377 8857 6411 8891
rect 6929 8857 6963 8891
rect 7849 8857 7883 8891
rect 10793 8857 10827 8891
rect 11989 8857 12023 8891
rect 13001 8857 13035 8891
rect 15209 8857 15243 8891
rect 17693 8857 17727 8891
rect 18107 8857 18141 8891
rect 2513 8789 2547 8823
rect 3433 8789 3467 8823
rect 5595 8789 5629 8823
rect 6469 8789 6503 8823
rect 8401 8789 8435 8823
rect 10885 8789 10919 8823
rect 16221 8789 16255 8823
rect 6101 8585 6135 8619
rect 8769 8585 8803 8619
rect 9413 8585 9447 8619
rect 13829 8585 13863 8619
rect 15853 8585 15887 8619
rect 9781 8517 9815 8551
rect 9919 8517 9953 8551
rect 12449 8517 12483 8551
rect 17969 8517 18003 8551
rect 2053 8449 2087 8483
rect 3617 8449 3651 8483
rect 4169 8449 4203 8483
rect 5733 8449 5767 8483
rect 6653 8449 6687 8483
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 7757 8449 7791 8483
rect 7941 8449 7975 8483
rect 8677 8449 8711 8483
rect 8861 8449 8895 8483
rect 9597 8449 9631 8483
rect 9689 8449 9723 8483
rect 10057 8449 10091 8483
rect 10517 8449 10551 8483
rect 10701 8449 10735 8483
rect 10793 8449 10827 8483
rect 11621 8449 11655 8483
rect 12357 8449 12391 8483
rect 12541 8449 12575 8483
rect 12817 8449 12851 8483
rect 13001 8449 13035 8483
rect 13645 8449 13679 8483
rect 13921 8449 13955 8483
rect 14197 8449 14231 8483
rect 14381 8449 14415 8483
rect 14657 8449 14691 8483
rect 14841 8449 14875 8483
rect 15485 8449 15519 8483
rect 16221 8449 16255 8483
rect 16808 8449 16842 8483
rect 2605 8381 2639 8415
rect 11713 8381 11747 8415
rect 12909 8381 12943 8415
rect 15853 8381 15887 8415
rect 4169 8313 4203 8347
rect 6101 8313 6135 8347
rect 6469 8313 6503 8347
rect 7113 8313 7147 8347
rect 13645 8313 13679 8347
rect 14289 8313 14323 8347
rect 18153 8313 18187 8347
rect 10333 8245 10367 8279
rect 14657 8245 14691 8279
rect 16313 8245 16347 8279
rect 16911 8245 16945 8279
rect 3433 8041 3467 8075
rect 6193 8041 6227 8075
rect 4721 7973 4755 8007
rect 7941 7973 7975 8007
rect 11345 7973 11379 8007
rect 12265 7973 12299 8007
rect 15301 7973 15335 8007
rect 3525 7905 3559 7939
rect 4261 7905 4295 7939
rect 4813 7905 4847 7939
rect 6009 7905 6043 7939
rect 6377 7905 6411 7939
rect 10333 7905 10367 7939
rect 11989 7905 12023 7939
rect 14289 7905 14323 7939
rect 14749 7905 14783 7939
rect 15577 7905 15611 7939
rect 2237 7837 2271 7871
rect 2329 7837 2363 7871
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 6745 7837 6779 7871
rect 7297 7837 7331 7871
rect 7665 7837 7699 7871
rect 7941 7837 7975 7871
rect 8125 7837 8159 7871
rect 10241 7837 10275 7871
rect 11253 7837 11287 7871
rect 11897 7837 11931 7871
rect 13277 7837 13311 7871
rect 13461 7837 13495 7871
rect 13579 7837 13613 7871
rect 13737 7837 13771 7871
rect 14381 7837 14415 7871
rect 15117 7837 15151 7871
rect 16497 7837 16531 7871
rect 16865 7837 16899 7871
rect 17785 7837 17819 7871
rect 18128 7837 18162 7871
rect 7389 7769 7423 7803
rect 13369 7769 13403 7803
rect 16221 7769 16255 7803
rect 17509 7769 17543 7803
rect 2053 7701 2087 7735
rect 6929 7701 6963 7735
rect 7481 7701 7515 7735
rect 7665 7701 7699 7735
rect 10609 7701 10643 7735
rect 13093 7701 13127 7735
rect 18199 7701 18233 7735
rect 5733 7497 5767 7531
rect 6863 7497 6897 7531
rect 8953 7497 8987 7531
rect 13369 7497 13403 7531
rect 16773 7497 16807 7531
rect 6653 7429 6687 7463
rect 15945 7429 15979 7463
rect 1685 7361 1719 7395
rect 1869 7361 1903 7395
rect 2421 7361 2455 7395
rect 2513 7361 2547 7395
rect 2605 7361 2639 7395
rect 2789 7361 2823 7395
rect 3249 7361 3283 7395
rect 4997 7361 5031 7395
rect 5641 7361 5675 7395
rect 5825 7361 5859 7395
rect 7665 7361 7699 7395
rect 7849 7361 7883 7395
rect 7941 7361 7975 7395
rect 8585 7361 8619 7395
rect 10333 7361 10367 7395
rect 11897 7361 11931 7395
rect 11989 7361 12023 7395
rect 12081 7361 12115 7395
rect 12265 7361 12299 7395
rect 13185 7361 13219 7395
rect 13921 7361 13955 7395
rect 15117 7361 15151 7395
rect 15301 7361 15335 7395
rect 15761 7361 15795 7395
rect 16957 7361 16991 7395
rect 17877 7361 17911 7395
rect 18153 7361 18187 7395
rect 1777 7293 1811 7327
rect 3065 7293 3099 7327
rect 4905 7293 4939 7327
rect 7757 7293 7791 7327
rect 8677 7293 8711 7327
rect 10425 7293 10459 7327
rect 11621 7293 11655 7327
rect 13001 7293 13035 7327
rect 13829 7293 13863 7327
rect 17233 7293 17267 7327
rect 5365 7225 5399 7259
rect 10701 7225 10735 7259
rect 14289 7225 14323 7259
rect 15117 7225 15151 7259
rect 2145 7157 2179 7191
rect 3433 7157 3467 7191
rect 6837 7157 6871 7191
rect 7021 7157 7055 7191
rect 7481 7157 7515 7191
rect 16129 7157 16163 7191
rect 4537 6953 4571 6987
rect 7941 6953 7975 6987
rect 7573 6885 7607 6919
rect 8125 6885 8159 6919
rect 9873 6885 9907 6919
rect 13461 6885 13495 6919
rect 2881 6817 2915 6851
rect 4261 6817 4295 6851
rect 6469 6817 6503 6851
rect 6745 6817 6779 6851
rect 10793 6817 10827 6851
rect 10977 6817 11011 6851
rect 11437 6817 11471 6851
rect 13001 6817 13035 6851
rect 14657 6817 14691 6851
rect 14841 6817 14875 6851
rect 16957 6817 16991 6851
rect 2421 6749 2455 6783
rect 2513 6749 2547 6783
rect 2605 6749 2639 6783
rect 4169 6749 4203 6783
rect 6377 6749 6411 6783
rect 8493 6749 8527 6783
rect 9502 6749 9536 6783
rect 9965 6749 9999 6783
rect 11529 6749 11563 6783
rect 12725 6749 12759 6783
rect 12817 6749 12851 6783
rect 13277 6749 13311 6783
rect 15209 6749 15243 6783
rect 15761 6749 15795 6783
rect 16405 6749 16439 6783
rect 16681 6749 16715 6783
rect 17233 6749 17267 6783
rect 18061 6749 18095 6783
rect 18429 6749 18463 6783
rect 2697 6681 2731 6715
rect 7941 6681 7975 6715
rect 8677 6681 8711 6715
rect 9321 6613 9355 6647
rect 9505 6613 9539 6647
rect 10333 6613 10367 6647
rect 10701 6613 10735 6647
rect 11897 6613 11931 6647
rect 13001 6613 13035 6647
rect 14197 6613 14231 6647
rect 14565 6613 14599 6647
rect 15393 6613 15427 6647
rect 18429 6613 18463 6647
rect 1869 6409 1903 6443
rect 2973 6409 3007 6443
rect 7849 6409 7883 6443
rect 9965 6409 9999 6443
rect 10977 6409 11011 6443
rect 14565 6409 14599 6443
rect 16313 6409 16347 6443
rect 2329 6341 2363 6375
rect 14473 6341 14507 6375
rect 15945 6341 15979 6375
rect 17693 6341 17727 6375
rect 2145 6273 2179 6307
rect 2237 6273 2271 6307
rect 3249 6273 3283 6307
rect 3341 6273 3375 6307
rect 3433 6273 3467 6307
rect 3617 6273 3651 6307
rect 3893 6273 3927 6307
rect 4077 6273 4111 6307
rect 4353 6273 4387 6307
rect 4537 6273 4571 6307
rect 4997 6273 5031 6307
rect 5181 6273 5215 6307
rect 5917 6273 5951 6307
rect 6101 6273 6135 6307
rect 6745 6273 6779 6307
rect 7757 6273 7791 6307
rect 8861 6273 8895 6307
rect 9597 6273 9631 6307
rect 9781 6273 9815 6307
rect 10425 6273 10459 6307
rect 10885 6273 10919 6307
rect 11621 6273 11655 6307
rect 12725 6273 12759 6307
rect 12817 6273 12851 6307
rect 13093 6273 13127 6307
rect 15761 6273 15795 6307
rect 16037 6273 16071 6307
rect 16129 6273 16163 6307
rect 17325 6273 17359 6307
rect 2605 6205 2639 6239
rect 6561 6205 6595 6239
rect 8033 6205 8067 6239
rect 9045 6205 9079 6239
rect 9137 6205 9171 6239
rect 13001 6205 13035 6239
rect 14749 6205 14783 6239
rect 10609 6137 10643 6171
rect 12541 6137 12575 6171
rect 17693 6137 17727 6171
rect 2513 6069 2547 6103
rect 5089 6069 5123 6103
rect 5917 6069 5951 6103
rect 6929 6069 6963 6103
rect 7389 6069 7423 6103
rect 8677 6069 8711 6103
rect 11805 6069 11839 6103
rect 13921 6069 13955 6103
rect 14105 6069 14139 6103
rect 2421 5865 2455 5899
rect 4169 5865 4203 5899
rect 4629 5865 4663 5899
rect 8585 5865 8619 5899
rect 9781 5865 9815 5899
rect 12909 5865 12943 5899
rect 13829 5865 13863 5899
rect 17969 5865 18003 5899
rect 4353 5797 4387 5831
rect 2789 5729 2823 5763
rect 4905 5729 4939 5763
rect 5089 5729 5123 5763
rect 7113 5729 7147 5763
rect 14197 5729 14231 5763
rect 14473 5729 14507 5763
rect 15945 5729 15979 5763
rect 16405 5729 16439 5763
rect 17049 5729 17083 5763
rect 1869 5661 1903 5695
rect 1961 5661 1995 5695
rect 2605 5661 2639 5695
rect 2697 5661 2731 5695
rect 2881 5661 2915 5695
rect 3065 5661 3099 5695
rect 4813 5661 4847 5695
rect 4997 5661 5031 5695
rect 5457 5661 5491 5695
rect 5611 5661 5645 5695
rect 6837 5661 6871 5695
rect 9321 5661 9355 5695
rect 9505 5661 9539 5695
rect 9781 5661 9815 5695
rect 9965 5661 9999 5695
rect 10333 5661 10367 5695
rect 11805 5661 11839 5695
rect 12633 5661 12667 5695
rect 12725 5661 12759 5695
rect 13185 5661 13219 5695
rect 13369 5661 13403 5695
rect 13645 5661 13679 5695
rect 17233 5661 17267 5695
rect 18153 5661 18187 5695
rect 3985 5593 4019 5627
rect 4201 5593 4235 5627
rect 10517 5593 10551 5627
rect 11897 5593 11931 5627
rect 13277 5593 13311 5627
rect 5825 5525 5859 5559
rect 8953 5525 8987 5559
rect 9413 5525 9447 5559
rect 2329 5321 2363 5355
rect 3249 5321 3283 5355
rect 4445 5321 4479 5355
rect 5365 5321 5399 5355
rect 6009 5321 6043 5355
rect 8033 5321 8067 5355
rect 8953 5321 8987 5355
rect 11069 5321 11103 5355
rect 13369 5321 13403 5355
rect 15485 5321 15519 5355
rect 16865 5321 16899 5355
rect 17233 5321 17267 5355
rect 1685 5253 1719 5287
rect 4721 5253 4755 5287
rect 9597 5253 9631 5287
rect 11897 5253 11931 5287
rect 14013 5253 14047 5287
rect 1593 5185 1627 5219
rect 2237 5185 2271 5219
rect 2421 5185 2455 5219
rect 3157 5185 3191 5219
rect 3341 5185 3375 5219
rect 4261 5185 4295 5219
rect 4905 5185 4939 5219
rect 4997 5185 5031 5219
rect 5273 5185 5307 5219
rect 5917 5185 5951 5219
rect 6101 5185 6135 5219
rect 6837 5185 6871 5219
rect 7941 5185 7975 5219
rect 8125 5185 8159 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 8861 5185 8895 5219
rect 9045 5185 9079 5219
rect 11621 5185 11655 5219
rect 13737 5185 13771 5219
rect 16037 5185 16071 5219
rect 16221 5185 16255 5219
rect 16773 5185 16807 5219
rect 16957 5185 16991 5219
rect 6929 5117 6963 5151
rect 7021 5117 7055 5151
rect 9321 5117 9355 5151
rect 4721 5049 4755 5083
rect 6469 4981 6503 5015
rect 8401 4981 8435 5015
rect 16037 4981 16071 5015
rect 7389 4777 7423 4811
rect 10793 4777 10827 4811
rect 11069 4777 11103 4811
rect 11345 4777 11379 4811
rect 11529 4777 11563 4811
rect 11713 4777 11747 4811
rect 12909 4777 12943 4811
rect 13645 4777 13679 4811
rect 13921 4777 13955 4811
rect 15945 4777 15979 4811
rect 3341 4641 3375 4675
rect 5917 4641 5951 4675
rect 8033 4641 8067 4675
rect 9321 4641 9355 4675
rect 14197 4641 14231 4675
rect 1685 4573 1719 4607
rect 1869 4573 1903 4607
rect 3249 4573 3283 4607
rect 4261 4573 4295 4607
rect 4813 4573 4847 4607
rect 5641 4573 5675 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 9045 4573 9079 4607
rect 11713 4573 11747 4607
rect 11897 4573 11931 4607
rect 12725 4573 12759 4607
rect 3157 4505 3191 4539
rect 12265 4505 12299 4539
rect 14473 4505 14507 4539
rect 2053 4437 2087 4471
rect 2789 4437 2823 4471
rect 4445 4437 4479 4471
rect 4997 4437 5031 4471
rect 7573 4437 7607 4471
rect 12357 4437 12391 4471
rect 4261 4233 4295 4267
rect 6653 4233 6687 4267
rect 11161 4233 11195 4267
rect 13645 4233 13679 4267
rect 2789 4165 2823 4199
rect 1685 4097 1719 4131
rect 1869 4097 1903 4131
rect 2053 4097 2087 4131
rect 2145 4097 2179 4131
rect 4537 4097 4571 4131
rect 4629 4097 4663 4131
rect 4721 4097 4755 4131
rect 5365 4097 5399 4131
rect 6561 4097 6595 4131
rect 6745 4097 6779 4131
rect 7205 4097 7239 4131
rect 9689 4097 9723 4131
rect 10149 4097 10183 4131
rect 10701 4097 10735 4131
rect 10885 4097 10919 4131
rect 11805 4097 11839 4131
rect 11989 4097 12023 4131
rect 13829 4097 13863 4131
rect 16129 4097 16163 4131
rect 16221 4097 16255 4131
rect 16313 4097 16347 4131
rect 17141 4097 17175 4131
rect 2513 4029 2547 4063
rect 4905 4029 4939 4063
rect 5457 4029 5491 4063
rect 7481 4029 7515 4063
rect 9229 4029 9263 4063
rect 9505 4029 9539 4063
rect 14105 4029 14139 4063
rect 17233 4029 17267 4063
rect 17417 4029 17451 4063
rect 16773 3961 16807 3995
rect 5641 3893 5675 3927
rect 9873 3893 9907 3927
rect 10333 3893 10367 3927
rect 10793 3893 10827 3927
rect 11805 3893 11839 3927
rect 15577 3893 15611 3927
rect 2789 3689 2823 3723
rect 5457 3689 5491 3723
rect 7665 3689 7699 3723
rect 8033 3689 8067 3723
rect 12173 3689 12207 3723
rect 13737 3689 13771 3723
rect 17049 3689 17083 3723
rect 5181 3621 5215 3655
rect 7205 3621 7239 3655
rect 17325 3621 17359 3655
rect 2145 3553 2179 3587
rect 2513 3553 2547 3587
rect 4721 3553 4755 3587
rect 8125 3553 8159 3587
rect 11897 3553 11931 3587
rect 14197 3553 14231 3587
rect 14473 3553 14507 3587
rect 17877 3553 17911 3587
rect 1685 3485 1719 3519
rect 2421 3485 2455 3519
rect 4859 3485 4893 3519
rect 5641 3485 5675 3519
rect 5733 3485 5767 3519
rect 5917 3485 5951 3519
rect 6009 3485 6043 3519
rect 6837 3485 6871 3519
rect 6991 3485 7025 3519
rect 7849 3485 7883 3519
rect 9505 3485 9539 3519
rect 9597 3485 9631 3519
rect 9689 3485 9723 3519
rect 9873 3485 9907 3519
rect 10149 3485 10183 3519
rect 13093 3485 13127 3519
rect 13277 3485 13311 3519
rect 16405 3485 16439 3519
rect 16773 3485 16807 3519
rect 16890 3485 16924 3519
rect 17785 3485 17819 3519
rect 2630 3417 2664 3451
rect 9229 3417 9263 3451
rect 10425 3417 10459 3451
rect 13185 3417 13219 3451
rect 13645 3417 13679 3451
rect 17693 3417 17727 3451
rect 1777 3349 1811 3383
rect 15945 3349 15979 3383
rect 16681 3349 16715 3383
rect 2605 3145 2639 3179
rect 3709 3145 3743 3179
rect 7021 3145 7055 3179
rect 8033 3145 8067 3179
rect 8861 3145 8895 3179
rect 9873 3145 9907 3179
rect 10977 3145 11011 3179
rect 13461 3145 13495 3179
rect 13737 3145 13771 3179
rect 15669 3145 15703 3179
rect 1777 3077 1811 3111
rect 5549 3077 5583 3111
rect 8493 3077 8527 3111
rect 8693 3077 8727 3111
rect 16313 3077 16347 3111
rect 1685 3009 1719 3043
rect 2237 3009 2271 3043
rect 2329 3009 2363 3043
rect 2421 3009 2455 3043
rect 3433 3009 3467 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 6653 3009 6687 3043
rect 6837 3009 6871 3043
rect 7481 3009 7515 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 9505 3009 9539 3043
rect 9659 3009 9693 3043
rect 10885 3009 10919 3043
rect 11713 3009 11747 3043
rect 13921 3009 13955 3043
rect 16221 3009 16255 3043
rect 16405 3009 16439 3043
rect 16957 3009 16991 3043
rect 17111 3009 17145 3043
rect 17693 3009 17727 3043
rect 3709 2941 3743 2975
rect 4997 2941 5031 2975
rect 11069 2941 11103 2975
rect 11989 2941 12023 2975
rect 14197 2941 14231 2975
rect 17325 2941 17359 2975
rect 10517 2873 10551 2907
rect 3525 2805 3559 2839
rect 4169 2805 4203 2839
rect 7481 2805 7515 2839
rect 8677 2805 8711 2839
rect 17785 2805 17819 2839
rect 1961 2601 1995 2635
rect 2605 2601 2639 2635
rect 3985 2601 4019 2635
rect 4537 2601 4571 2635
rect 5825 2601 5859 2635
rect 6377 2601 6411 2635
rect 11621 2601 11655 2635
rect 13001 2601 13035 2635
rect 3433 2533 3467 2567
rect 7849 2533 7883 2567
rect 9137 2533 9171 2567
rect 16037 2533 16071 2567
rect 9321 2465 9355 2499
rect 15761 2465 15795 2499
rect 1777 2397 1811 2431
rect 1870 2397 1904 2431
rect 2605 2397 2639 2431
rect 2789 2397 2823 2431
rect 3157 2397 3191 2431
rect 3249 2397 3283 2431
rect 3893 2397 3927 2431
rect 4077 2397 4111 2431
rect 4537 2397 4571 2431
rect 4813 2397 4847 2431
rect 5457 2397 5491 2431
rect 5641 2397 5675 2431
rect 6377 2397 6411 2431
rect 6561 2397 6595 2431
rect 6929 2397 6963 2431
rect 7113 2397 7147 2431
rect 8125 2397 8159 2431
rect 8677 2397 8711 2431
rect 9045 2397 9079 2431
rect 9873 2397 9907 2431
rect 13001 2397 13035 2431
rect 13185 2397 13219 2431
rect 14197 2397 14231 2431
rect 14381 2397 14415 2431
rect 14841 2397 14875 2431
rect 15025 2397 15059 2431
rect 15669 2397 15703 2431
rect 7849 2329 7883 2363
rect 8033 2329 8067 2363
rect 8493 2329 8527 2363
rect 10149 2329 10183 2363
rect 4721 2261 4755 2295
rect 7021 2261 7055 2295
rect 9321 2261 9355 2295
rect 11805 2261 11839 2295
rect 11989 2261 12023 2295
rect 13737 2261 13771 2295
rect 14289 2261 14323 2295
rect 14933 2261 14967 2295
rect 3709 2057 3743 2091
rect 6101 2057 6135 2091
rect 10885 2057 10919 2091
rect 13461 2057 13495 2091
rect 6469 1989 6503 2023
rect 14013 1989 14047 2023
rect 1961 1921 1995 1955
rect 4077 1921 4111 1955
rect 6653 1921 6687 1955
rect 6745 1921 6779 1955
rect 7665 1921 7699 1955
rect 8401 1921 8435 1955
rect 10793 1921 10827 1955
rect 10977 1921 11011 1955
rect 2237 1853 2271 1887
rect 4353 1853 4387 1887
rect 7573 1853 7607 1887
rect 8677 1853 8711 1887
rect 10425 1853 10459 1887
rect 11713 1853 11747 1887
rect 11989 1853 12023 1887
rect 13737 1853 13771 1887
rect 5825 1785 5859 1819
rect 6561 1717 6595 1751
rect 7941 1717 7975 1751
rect 11253 1717 11287 1751
rect 15485 1717 15519 1751
rect 2329 1513 2363 1547
rect 3893 1513 3927 1547
rect 4261 1513 4295 1547
rect 4905 1513 4939 1547
rect 6726 1513 6760 1547
rect 8217 1513 8251 1547
rect 8401 1513 8435 1547
rect 9505 1513 9539 1547
rect 10701 1513 10735 1547
rect 13553 1513 13587 1547
rect 13829 1513 13863 1547
rect 15945 1513 15979 1547
rect 2605 1445 2639 1479
rect 10517 1445 10551 1479
rect 10977 1445 11011 1479
rect 11897 1445 11931 1479
rect 3249 1377 3283 1411
rect 5457 1377 5491 1411
rect 6469 1377 6503 1411
rect 14197 1377 14231 1411
rect 14473 1377 14507 1411
rect 1777 1309 1811 1343
rect 2973 1309 3007 1343
rect 3065 1309 3099 1343
rect 4261 1309 4295 1343
rect 4445 1309 4479 1343
rect 5273 1309 5307 1343
rect 9321 1309 9355 1343
rect 9781 1309 9815 1343
rect 10241 1309 10275 1343
rect 10333 1309 10367 1343
rect 10977 1309 11011 1343
rect 11161 1309 11195 1343
rect 11897 1309 11931 1343
rect 12081 1309 12115 1343
rect 5365 1241 5399 1275
rect 1961 1173 1995 1207
rect 9689 1173 9723 1207
<< metal1 >>
rect 1394 14288 1400 14340
rect 1452 14328 1458 14340
rect 7098 14328 7104 14340
rect 1452 14300 7104 14328
rect 1452 14288 1458 14300
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 1104 13626 18860 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 18860 13626
rect 1104 13552 18860 13574
rect 12250 13512 12256 13524
rect 3896 13484 12256 13512
rect 3050 13336 3056 13388
rect 3108 13376 3114 13388
rect 3896 13385 3924 13484
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 4249 13447 4307 13453
rect 4249 13413 4261 13447
rect 4295 13444 4307 13447
rect 4709 13447 4767 13453
rect 4709 13444 4721 13447
rect 4295 13416 4721 13444
rect 4295 13413 4307 13416
rect 4249 13407 4307 13413
rect 4709 13413 4721 13416
rect 4755 13413 4767 13447
rect 4709 13407 4767 13413
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 9033 13447 9091 13453
rect 9033 13444 9045 13447
rect 8527 13416 9045 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9033 13413 9045 13416
rect 9079 13413 9091 13447
rect 9033 13407 9091 13413
rect 13081 13447 13139 13453
rect 13081 13413 13093 13447
rect 13127 13444 13139 13447
rect 13357 13447 13415 13453
rect 13357 13444 13369 13447
rect 13127 13416 13369 13444
rect 13127 13413 13139 13416
rect 13081 13407 13139 13413
rect 13357 13413 13369 13416
rect 13403 13413 13415 13447
rect 13357 13407 13415 13413
rect 16347 13447 16405 13453
rect 16347 13413 16359 13447
rect 16393 13444 16405 13447
rect 16393 13416 16574 13444
rect 16393 13413 16405 13416
rect 16347 13407 16405 13413
rect 3881 13379 3939 13385
rect 3881 13376 3893 13379
rect 3108 13348 3893 13376
rect 3108 13336 3114 13348
rect 3881 13345 3893 13348
rect 3927 13345 3939 13379
rect 3881 13339 3939 13345
rect 6549 13379 6607 13385
rect 6549 13345 6561 13379
rect 6595 13376 6607 13379
rect 6914 13376 6920 13388
rect 6595 13348 6920 13376
rect 6595 13345 6607 13348
rect 6549 13339 6607 13345
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 7834 13336 7840 13388
rect 7892 13376 7898 13388
rect 9631 13379 9689 13385
rect 9631 13376 9643 13379
rect 7892 13348 9643 13376
rect 7892 13336 7898 13348
rect 9631 13345 9643 13348
rect 9677 13345 9689 13379
rect 16546 13376 16574 13416
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 9631 13339 9689 13345
rect 9784 13348 15608 13376
rect 16546 13348 17325 13376
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4120 13280 4905 13308
rect 4120 13268 4126 13280
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5691 13311 5749 13317
rect 5691 13277 5703 13311
rect 5737 13308 5749 13311
rect 5737 13280 5856 13308
rect 5737 13277 5749 13280
rect 5691 13271 5749 13277
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13172 4307 13175
rect 4798 13172 4804 13184
rect 4295 13144 4804 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 5828 13172 5856 13280
rect 6730 13268 6736 13320
rect 6788 13268 6794 13320
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7098 13308 7104 13320
rect 7055 13280 7104 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 8110 13268 8116 13320
rect 8168 13268 8174 13320
rect 9214 13268 9220 13320
rect 9272 13268 9278 13320
rect 9528 13311 9586 13317
rect 9528 13308 9540 13311
rect 9324 13280 9540 13308
rect 5905 13243 5963 13249
rect 5905 13209 5917 13243
rect 5951 13240 5963 13243
rect 7282 13240 7288 13252
rect 5951 13212 7288 13240
rect 5951 13209 5963 13212
rect 5905 13203 5963 13209
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 7377 13243 7435 13249
rect 7377 13209 7389 13243
rect 7423 13240 7435 13243
rect 9122 13240 9128 13252
rect 7423 13212 9128 13240
rect 7423 13209 7435 13212
rect 7377 13203 7435 13209
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 6917 13175 6975 13181
rect 6917 13172 6929 13175
rect 5828 13144 6929 13172
rect 6917 13141 6929 13144
rect 6963 13172 6975 13175
rect 7190 13172 7196 13184
rect 6963 13144 7196 13172
rect 6963 13141 6975 13144
rect 6917 13135 6975 13141
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 7466 13132 7472 13184
rect 7524 13132 7530 13184
rect 8481 13175 8539 13181
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 8662 13172 8668 13184
rect 8527 13144 8668 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 8662 13132 8668 13144
rect 8720 13172 8726 13184
rect 9324 13172 9352 13280
rect 9528 13277 9540 13280
rect 9574 13277 9586 13311
rect 9528 13271 9586 13277
rect 9398 13200 9404 13252
rect 9456 13240 9462 13252
rect 9784 13240 9812 13348
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 9456 13212 9812 13240
rect 10244 13240 10272 13271
rect 10318 13268 10324 13320
rect 10376 13268 10382 13320
rect 12044 13311 12102 13317
rect 12044 13277 12056 13311
rect 12090 13308 12102 13311
rect 12090 13280 12664 13308
rect 12090 13277 12102 13280
rect 12044 13271 12102 13277
rect 10410 13240 10416 13252
rect 10244 13212 10416 13240
rect 9456 13200 9462 13212
rect 10410 13200 10416 13212
rect 10468 13200 10474 13252
rect 8720 13144 9352 13172
rect 8720 13132 8726 13144
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10229 13175 10287 13181
rect 10229 13172 10241 13175
rect 10100 13144 10241 13172
rect 10100 13132 10106 13144
rect 10229 13141 10241 13144
rect 10275 13172 10287 13175
rect 10594 13172 10600 13184
rect 10275 13144 10600 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 12158 13181 12164 13184
rect 12115 13175 12164 13181
rect 12115 13141 12127 13175
rect 12161 13141 12164 13175
rect 12115 13135 12164 13141
rect 12158 13132 12164 13135
rect 12216 13132 12222 13184
rect 12636 13172 12664 13280
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 13541 13311 13599 13317
rect 13541 13308 13553 13311
rect 13504 13280 13553 13308
rect 13504 13268 13510 13280
rect 13541 13277 13553 13280
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 14185 13311 14243 13317
rect 14185 13277 14197 13311
rect 14231 13308 14243 13311
rect 14458 13308 14464 13320
rect 14231 13280 14464 13308
rect 14231 13277 14243 13280
rect 14185 13271 14243 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 15580 13317 15608 13348
rect 17313 13345 17325 13348
rect 17359 13345 17371 13379
rect 17313 13339 17371 13345
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 16276 13311 16334 13317
rect 16276 13277 16288 13311
rect 16322 13308 16334 13311
rect 16666 13308 16672 13320
rect 16322 13280 16672 13308
rect 16322 13277 16334 13280
rect 16276 13271 16334 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 16758 13268 16764 13320
rect 16816 13268 16822 13320
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 17144 13280 17785 13308
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 14645 13243 14703 13249
rect 14645 13240 14657 13243
rect 14608 13212 14657 13240
rect 14608 13200 14614 13212
rect 14645 13209 14657 13212
rect 14691 13209 14703 13243
rect 14645 13203 14703 13209
rect 14734 13200 14740 13252
rect 14792 13200 14798 13252
rect 15749 13243 15807 13249
rect 15749 13209 15761 13243
rect 15795 13240 15807 13243
rect 16114 13240 16120 13252
rect 15795 13212 16120 13240
rect 15795 13209 15807 13212
rect 15749 13203 15807 13209
rect 16114 13200 16120 13212
rect 16172 13240 16178 13252
rect 17144 13240 17172 13280
rect 17773 13277 17785 13280
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 16172 13212 17172 13240
rect 17221 13243 17279 13249
rect 16172 13200 16178 13212
rect 17221 13209 17233 13243
rect 17267 13240 17279 13243
rect 17402 13240 17408 13252
rect 17267 13212 17408 13240
rect 17267 13209 17279 13212
rect 17221 13203 17279 13209
rect 17402 13200 17408 13212
rect 17460 13200 17466 13252
rect 13081 13175 13139 13181
rect 13081 13172 13093 13175
rect 12636 13144 13093 13172
rect 13081 13141 13093 13144
rect 13127 13172 13139 13175
rect 13354 13172 13360 13184
rect 13127 13144 13360 13172
rect 13127 13141 13139 13144
rect 13081 13135 13139 13141
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 15286 13172 15292 13184
rect 13688 13144 15292 13172
rect 13688 13132 13694 13144
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 17586 13132 17592 13184
rect 17644 13132 17650 13184
rect 1104 13082 18860 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 16214 13082
rect 16266 13030 16278 13082
rect 16330 13030 16342 13082
rect 16394 13030 16406 13082
rect 16458 13030 16470 13082
rect 16522 13030 18860 13082
rect 1104 13008 18860 13030
rect 8662 12928 8668 12980
rect 8720 12928 8726 12980
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 11054 12968 11060 12980
rect 9180 12940 11060 12968
rect 9180 12928 9186 12940
rect 11054 12928 11060 12940
rect 11112 12968 11118 12980
rect 11112 12940 12112 12968
rect 11112 12928 11118 12940
rect 4341 12903 4399 12909
rect 4341 12869 4353 12903
rect 4387 12900 4399 12903
rect 4614 12900 4620 12912
rect 4387 12872 4620 12900
rect 4387 12869 4399 12872
rect 4341 12863 4399 12869
rect 4614 12860 4620 12872
rect 4672 12900 4678 12912
rect 5813 12903 5871 12909
rect 5813 12900 5825 12903
rect 4672 12872 5825 12900
rect 4672 12860 4678 12872
rect 5813 12869 5825 12872
rect 5859 12869 5871 12903
rect 5813 12863 5871 12869
rect 7742 12860 7748 12912
rect 7800 12900 7806 12912
rect 9398 12900 9404 12912
rect 7800 12872 9404 12900
rect 7800 12860 7806 12872
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 9999 12903 10057 12909
rect 9999 12869 10011 12903
rect 10045 12900 10057 12903
rect 10134 12900 10140 12912
rect 10045 12872 10140 12900
rect 10045 12869 10057 12872
rect 9999 12863 10057 12869
rect 10134 12860 10140 12872
rect 10192 12860 10198 12912
rect 12084 12909 12112 12940
rect 12250 12928 12256 12980
rect 12308 12968 12314 12980
rect 13170 12968 13176 12980
rect 12308 12940 13176 12968
rect 12308 12928 12314 12940
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 13354 12928 13360 12980
rect 13412 12928 13418 12980
rect 15470 12928 15476 12980
rect 15528 12968 15534 12980
rect 16758 12968 16764 12980
rect 15528 12940 16764 12968
rect 15528 12928 15534 12940
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 10689 12903 10747 12909
rect 10689 12900 10701 12903
rect 10612 12872 10701 12900
rect 10612 12844 10640 12872
rect 10689 12869 10701 12872
rect 10735 12869 10747 12903
rect 10689 12863 10747 12869
rect 12069 12903 12127 12909
rect 12069 12869 12081 12903
rect 12115 12869 12127 12903
rect 12069 12863 12127 12869
rect 12158 12860 12164 12912
rect 12216 12860 12222 12912
rect 14366 12860 14372 12912
rect 14424 12900 14430 12912
rect 14424 12872 16068 12900
rect 14424 12860 14430 12872
rect 3050 12792 3056 12844
rect 3108 12792 3114 12844
rect 3602 12792 3608 12844
rect 3660 12792 3666 12844
rect 3878 12792 3884 12844
rect 3936 12792 3942 12844
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12832 6515 12835
rect 6914 12832 6920 12844
rect 6503 12804 6920 12832
rect 6503 12801 6515 12804
rect 6457 12795 6515 12801
rect 3620 12764 3648 12792
rect 4062 12764 4068 12776
rect 3620 12736 4068 12764
rect 4062 12724 4068 12736
rect 4120 12764 4126 12776
rect 4448 12764 4476 12795
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 4120 12736 4476 12764
rect 5997 12767 6055 12773
rect 4120 12724 4126 12736
rect 5997 12733 6009 12767
rect 6043 12764 6055 12767
rect 7024 12764 7052 12795
rect 8110 12792 8116 12844
rect 8168 12832 8174 12844
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 8168 12804 8309 12832
rect 8168 12792 8174 12804
rect 8297 12801 8309 12804
rect 8343 12832 8355 12835
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 8343 12804 9505 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 9493 12801 9505 12804
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 9674 12792 9680 12844
rect 9732 12792 9738 12844
rect 9766 12792 9772 12844
rect 9824 12792 9830 12844
rect 9858 12792 9864 12844
rect 9916 12792 9922 12844
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10505 12835 10563 12841
rect 10505 12832 10517 12835
rect 10284 12804 10517 12832
rect 10284 12792 10290 12804
rect 10505 12801 10517 12804
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 10594 12792 10600 12844
rect 10652 12792 10658 12844
rect 10962 12841 10968 12844
rect 10773 12835 10831 12841
rect 10773 12832 10785 12835
rect 10704 12804 10785 12832
rect 8665 12767 8723 12773
rect 8665 12764 8677 12767
rect 6043 12736 8677 12764
rect 6043 12733 6055 12736
rect 5997 12727 6055 12733
rect 8665 12733 8677 12736
rect 8711 12764 8723 12767
rect 9214 12764 9220 12776
rect 8711 12736 9220 12764
rect 8711 12733 8723 12736
rect 8665 12727 8723 12733
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 10410 12764 10416 12776
rect 10183 12736 10416 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10410 12724 10416 12736
rect 10468 12764 10474 12776
rect 10704 12764 10732 12804
rect 10773 12801 10785 12804
rect 10819 12801 10831 12835
rect 10773 12795 10831 12801
rect 10919 12835 10968 12841
rect 10919 12801 10931 12835
rect 10965 12801 10968 12835
rect 10919 12795 10968 12801
rect 10962 12792 10968 12795
rect 11020 12792 11026 12844
rect 14458 12792 14464 12844
rect 14516 12832 14522 12844
rect 14645 12835 14703 12841
rect 14645 12832 14657 12835
rect 14516 12804 14657 12832
rect 14516 12792 14522 12804
rect 14645 12801 14657 12804
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 15194 12792 15200 12844
rect 15252 12792 15258 12844
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 15344 12804 15761 12832
rect 15344 12792 15350 12804
rect 15749 12801 15761 12804
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 15930 12792 15936 12844
rect 15988 12792 15994 12844
rect 16040 12841 16068 12872
rect 16666 12860 16672 12912
rect 16724 12900 16730 12912
rect 17221 12903 17279 12909
rect 17221 12900 17233 12903
rect 16724 12872 17233 12900
rect 16724 12860 16730 12872
rect 17221 12869 17233 12872
rect 17267 12900 17279 12903
rect 17678 12900 17684 12912
rect 17267 12872 17684 12900
rect 17267 12869 17279 12872
rect 17221 12863 17279 12869
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 16758 12792 16764 12844
rect 16816 12792 16822 12844
rect 18046 12841 18052 12844
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12801 17371 12835
rect 17313 12795 17371 12801
rect 18024 12835 18052 12841
rect 18024 12801 18036 12835
rect 18024 12795 18052 12801
rect 10468 12736 10732 12764
rect 10468 12724 10474 12736
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 11204 12736 11621 12764
rect 11204 12724 11210 12736
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 12710 12724 12716 12776
rect 12768 12764 12774 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12768 12736 13001 12764
rect 12768 12724 12774 12736
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 3605 12699 3663 12705
rect 3605 12665 3617 12699
rect 3651 12696 3663 12699
rect 4798 12696 4804 12708
rect 3651 12668 4804 12696
rect 3651 12665 3663 12668
rect 3605 12659 3663 12665
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 7009 12699 7067 12705
rect 7009 12665 7021 12699
rect 7055 12696 7067 12699
rect 7742 12696 7748 12708
rect 7055 12668 7748 12696
rect 7055 12665 7067 12668
rect 7009 12659 7067 12665
rect 7742 12656 7748 12668
rect 7800 12656 7806 12708
rect 13004 12696 13032 12727
rect 13354 12724 13360 12776
rect 13412 12724 13418 12776
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14550 12764 14556 12776
rect 14148 12736 14556 12764
rect 14148 12724 14154 12736
rect 14550 12724 14556 12736
rect 14608 12764 14614 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14608 12736 15025 12764
rect 14608 12724 14614 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 16114 12724 16120 12776
rect 16172 12764 16178 12776
rect 17328 12764 17356 12795
rect 18046 12792 18052 12795
rect 18104 12792 18110 12844
rect 16172 12736 17356 12764
rect 16172 12724 16178 12736
rect 15565 12699 15623 12705
rect 15565 12696 15577 12699
rect 13004 12668 15577 12696
rect 15565 12665 15577 12668
rect 15611 12665 15623 12699
rect 15565 12659 15623 12665
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 15470 12628 15476 12640
rect 11103 12600 15476 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 18095 12631 18153 12637
rect 18095 12597 18107 12631
rect 18141 12628 18153 12631
rect 18230 12628 18236 12640
rect 18141 12600 18236 12628
rect 18141 12597 18153 12600
rect 18095 12591 18153 12597
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 1104 12538 18860 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 18860 12538
rect 1104 12464 18860 12486
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 9858 12424 9864 12436
rect 3292 12396 9864 12424
rect 3292 12384 3298 12396
rect 9858 12384 9864 12396
rect 9916 12424 9922 12436
rect 9953 12427 10011 12433
rect 9953 12424 9965 12427
rect 9916 12396 9965 12424
rect 9916 12384 9922 12396
rect 9953 12393 9965 12396
rect 9999 12393 10011 12427
rect 13078 12424 13084 12436
rect 9953 12387 10011 12393
rect 10060 12396 13084 12424
rect 2685 12359 2743 12365
rect 2685 12325 2697 12359
rect 2731 12356 2743 12359
rect 2866 12356 2872 12368
rect 2731 12328 2872 12356
rect 2731 12325 2743 12328
rect 2685 12319 2743 12325
rect 2866 12316 2872 12328
rect 2924 12316 2930 12368
rect 3142 12316 3148 12368
rect 3200 12356 3206 12368
rect 3602 12356 3608 12368
rect 3200 12328 3608 12356
rect 3200 12316 3206 12328
rect 3602 12316 3608 12328
rect 3660 12316 3666 12368
rect 4614 12316 4620 12368
rect 4672 12316 4678 12368
rect 7742 12316 7748 12368
rect 7800 12316 7806 12368
rect 7926 12316 7932 12368
rect 7984 12356 7990 12368
rect 10060 12356 10088 12396
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13170 12384 13176 12436
rect 13228 12384 13234 12436
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13412 12396 13737 12424
rect 13412 12384 13418 12396
rect 13725 12393 13737 12396
rect 13771 12393 13783 12427
rect 13725 12387 13783 12393
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 15151 12427 15209 12433
rect 15151 12424 15163 12427
rect 14792 12396 15163 12424
rect 14792 12384 14798 12396
rect 15151 12393 15163 12396
rect 15197 12393 15209 12427
rect 15151 12387 15209 12393
rect 16025 12427 16083 12433
rect 16025 12393 16037 12427
rect 16071 12424 16083 12427
rect 17402 12424 17408 12436
rect 16071 12396 17408 12424
rect 16071 12393 16083 12396
rect 16025 12387 16083 12393
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 17678 12384 17684 12436
rect 17736 12384 17742 12436
rect 13372 12356 13400 12384
rect 18782 12356 18788 12368
rect 7984 12328 10088 12356
rect 11256 12328 13400 12356
rect 13556 12328 18788 12356
rect 7984 12316 7990 12328
rect 3053 12291 3111 12297
rect 1872 12260 3004 12288
rect 1872 12229 1900 12260
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12189 1915 12223
rect 1857 12183 1915 12189
rect 2130 12180 2136 12232
rect 2188 12180 2194 12232
rect 2222 12112 2228 12164
rect 2280 12152 2286 12164
rect 2501 12155 2559 12161
rect 2501 12152 2513 12155
rect 2280 12124 2513 12152
rect 2280 12112 2286 12124
rect 2501 12121 2513 12124
rect 2547 12121 2559 12155
rect 2976 12152 3004 12260
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 3878 12288 3884 12300
rect 3099 12260 3884 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 3878 12248 3884 12260
rect 3936 12288 3942 12300
rect 4157 12291 4215 12297
rect 4157 12288 4169 12291
rect 3936 12260 4169 12288
rect 3936 12248 3942 12260
rect 4157 12257 4169 12260
rect 4203 12257 4215 12291
rect 4157 12251 4215 12257
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 6972 12260 7297 12288
rect 6972 12248 6978 12260
rect 7285 12257 7297 12260
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 7834 12248 7840 12300
rect 7892 12248 7898 12300
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12288 8263 12291
rect 8251 12260 10732 12288
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3510 12180 3516 12232
rect 3568 12180 3574 12232
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 5020 12223 5078 12229
rect 5020 12220 5032 12223
rect 4856 12192 5032 12220
rect 4856 12180 4862 12192
rect 5020 12189 5032 12192
rect 5066 12189 5078 12223
rect 5020 12183 5078 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 3878 12152 3884 12164
rect 2976 12124 3884 12152
rect 2501 12115 2559 12121
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 4709 12155 4767 12161
rect 4709 12121 4721 12155
rect 4755 12152 4767 12155
rect 5123 12155 5181 12161
rect 5123 12152 5135 12155
rect 4755 12124 5135 12152
rect 4755 12121 4767 12124
rect 4709 12115 4767 12121
rect 5123 12121 5135 12124
rect 5169 12121 5181 12155
rect 6288 12152 6316 12183
rect 6638 12180 6644 12232
rect 6696 12180 6702 12232
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12220 8723 12223
rect 8846 12220 8852 12232
rect 8711 12192 8852 12220
rect 8711 12189 8723 12192
rect 8665 12183 8723 12189
rect 7926 12152 7932 12164
rect 6288 12124 7932 12152
rect 5123 12115 5181 12121
rect 7926 12112 7932 12124
rect 7984 12112 7990 12164
rect 8404 12152 8432 12183
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 10134 12220 10140 12232
rect 9447 12192 10140 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12220 10287 12223
rect 10318 12220 10324 12232
rect 10275 12192 10324 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10704 12229 10732 12260
rect 11054 12248 11060 12300
rect 11112 12248 11118 12300
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12220 10747 12223
rect 11146 12220 11152 12232
rect 10735 12192 11152 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11256 12229 11284 12328
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 11572 12192 12173 12220
rect 11572 12180 11578 12192
rect 12161 12189 12173 12192
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13556 12220 13584 12328
rect 18782 12316 18788 12328
rect 18840 12316 18846 12368
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 17644 12260 17693 12288
rect 17644 12248 17650 12260
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 17681 12251 17739 12257
rect 13035 12192 13584 12220
rect 13633 12223 13691 12229
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13633 12189 13645 12223
rect 13679 12220 13691 12223
rect 14090 12220 14096 12232
rect 13679 12192 14096 12220
rect 13679 12189 13691 12192
rect 13633 12183 13691 12189
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14182 12180 14188 12232
rect 14240 12180 14246 12232
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12220 14611 12223
rect 14826 12220 14832 12232
rect 14599 12192 14832 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15048 12223 15106 12229
rect 15048 12220 15060 12223
rect 14936 12192 15060 12220
rect 9953 12155 10011 12161
rect 8404 12124 8708 12152
rect 8680 12096 8708 12124
rect 9953 12121 9965 12155
rect 9999 12152 10011 12155
rect 10410 12152 10416 12164
rect 9999 12124 10416 12152
rect 9999 12121 10011 12124
rect 9953 12115 10011 12121
rect 10410 12112 10416 12124
rect 10468 12152 10474 12164
rect 10778 12152 10784 12164
rect 10468 12124 10784 12152
rect 10468 12112 10474 12124
rect 10778 12112 10784 12124
rect 10836 12112 10842 12164
rect 11790 12112 11796 12164
rect 11848 12152 11854 12164
rect 12805 12155 12863 12161
rect 12805 12152 12817 12155
rect 11848 12124 12817 12152
rect 11848 12112 11854 12124
rect 12805 12121 12817 12124
rect 12851 12121 12863 12155
rect 12805 12115 12863 12121
rect 12897 12155 12955 12161
rect 12897 12121 12909 12155
rect 12943 12152 12955 12155
rect 14366 12152 14372 12164
rect 12943 12124 14372 12152
rect 12943 12121 12955 12124
rect 12897 12115 12955 12121
rect 14366 12112 14372 12124
rect 14424 12112 14430 12164
rect 14936 12152 14964 12192
rect 15048 12189 15060 12192
rect 15094 12189 15106 12223
rect 15048 12183 15106 12189
rect 15470 12180 15476 12232
rect 15528 12180 15534 12232
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12220 16083 12223
rect 16114 12220 16120 12232
rect 16071 12192 16120 12220
rect 16071 12189 16083 12192
rect 16025 12183 16083 12189
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 17310 12220 17316 12232
rect 16816 12192 17316 12220
rect 16816 12180 16822 12192
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 17460 12192 18245 12220
rect 17460 12180 17466 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 14568 12124 14964 12152
rect 14568 12096 14596 12124
rect 1486 12044 1492 12096
rect 1544 12084 1550 12096
rect 1673 12087 1731 12093
rect 1673 12084 1685 12087
rect 1544 12056 1685 12084
rect 1544 12044 1550 12056
rect 1673 12053 1685 12056
rect 1719 12053 1731 12087
rect 1673 12047 1731 12053
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 2130 12084 2136 12096
rect 2087 12056 2136 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 2130 12044 2136 12056
rect 2188 12084 2194 12096
rect 3418 12084 3424 12096
rect 2188 12056 3424 12084
rect 2188 12044 2194 12056
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 6641 12087 6699 12093
rect 6641 12084 6653 12087
rect 6604 12056 6653 12084
rect 6604 12044 6610 12056
rect 6641 12053 6653 12056
rect 6687 12053 6699 12087
rect 6641 12047 6699 12053
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 8076 12056 8585 12084
rect 8076 12044 8082 12056
rect 8573 12053 8585 12056
rect 8619 12053 8631 12087
rect 8573 12047 8631 12053
rect 8662 12044 8668 12096
rect 8720 12044 8726 12096
rect 9306 12044 9312 12096
rect 9364 12044 9370 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 10137 12087 10195 12093
rect 10137 12084 10149 12087
rect 9456 12056 10149 12084
rect 9456 12044 9462 12056
rect 10137 12053 10149 12056
rect 10183 12053 10195 12087
rect 10137 12047 10195 12053
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 11146 12084 11152 12096
rect 10376 12056 11152 12084
rect 10376 12044 10382 12056
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 12710 12084 12716 12096
rect 12391 12056 12716 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 14550 12044 14556 12096
rect 14608 12044 14614 12096
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 18325 12087 18383 12093
rect 18325 12084 18337 12087
rect 17460 12056 18337 12084
rect 17460 12044 17466 12056
rect 18325 12053 18337 12056
rect 18371 12053 18383 12087
rect 18325 12047 18383 12053
rect 1104 11994 18860 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 16214 11994
rect 16266 11942 16278 11994
rect 16330 11942 16342 11994
rect 16394 11942 16406 11994
rect 16458 11942 16470 11994
rect 16522 11942 18860 11994
rect 1104 11920 18860 11942
rect 3418 11840 3424 11892
rect 3476 11880 3482 11892
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 3476 11852 4629 11880
rect 3476 11840 3482 11852
rect 4617 11849 4629 11852
rect 4663 11849 4675 11883
rect 4617 11843 4675 11849
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 6638 11880 6644 11892
rect 5951 11852 6644 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 8018 11880 8024 11892
rect 7248 11852 8024 11880
rect 7248 11840 7254 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 10042 11880 10048 11892
rect 8680 11852 10048 11880
rect 3694 11772 3700 11824
rect 3752 11812 3758 11824
rect 8481 11815 8539 11821
rect 8481 11812 8493 11815
rect 3752 11784 4752 11812
rect 3752 11772 3758 11784
rect 1486 11704 1492 11756
rect 1544 11704 1550 11756
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11744 2099 11747
rect 3510 11744 3516 11756
rect 2087 11716 3516 11744
rect 2087 11713 2099 11716
rect 2041 11707 2099 11713
rect 3510 11704 3516 11716
rect 3568 11744 3574 11756
rect 4433 11747 4491 11753
rect 3568 11716 3648 11744
rect 3568 11704 3574 11716
rect 3620 11676 3648 11716
rect 4433 11713 4445 11747
rect 4479 11744 4491 11747
rect 4614 11744 4620 11756
rect 4479 11716 4620 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 4724 11753 4752 11784
rect 7852 11784 8493 11812
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 5074 11704 5080 11756
rect 5132 11704 5138 11756
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5868 11716 6101 11744
rect 5868 11704 5874 11716
rect 6089 11713 6101 11716
rect 6135 11744 6147 11747
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 6135 11716 7389 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 7377 11713 7389 11716
rect 7423 11744 7435 11747
rect 7466 11744 7472 11756
rect 7423 11716 7472 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 7852 11753 7880 11784
rect 8481 11781 8493 11784
rect 8527 11781 8539 11815
rect 8481 11775 8539 11781
rect 8680 11756 8708 11852
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10962 11880 10968 11892
rect 10376 11852 10968 11880
rect 10376 11840 10382 11852
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 12805 11883 12863 11889
rect 12805 11849 12817 11883
rect 12851 11880 12863 11883
rect 14001 11883 14059 11889
rect 12851 11852 13676 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 11882 11812 11888 11824
rect 8812 11784 11888 11812
rect 8812 11772 8818 11784
rect 11882 11772 11888 11784
rect 11940 11772 11946 11824
rect 12437 11815 12495 11821
rect 12437 11781 12449 11815
rect 12483 11812 12495 11815
rect 13446 11812 13452 11824
rect 12483 11784 13452 11812
rect 12483 11781 12495 11784
rect 12437 11775 12495 11781
rect 13446 11772 13452 11784
rect 13504 11772 13510 11824
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 8570 11744 8576 11756
rect 8159 11716 8576 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8570 11704 8576 11716
rect 8628 11704 8634 11756
rect 8662 11704 8668 11756
rect 8720 11704 8726 11756
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11744 8907 11747
rect 9030 11744 9036 11756
rect 8895 11716 9036 11744
rect 8895 11713 8907 11716
rect 8849 11707 8907 11713
rect 5261 11679 5319 11685
rect 5261 11676 5273 11679
rect 3620 11648 5273 11676
rect 5261 11645 5273 11648
rect 5307 11645 5319 11679
rect 5261 11639 5319 11645
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 7926 11676 7932 11688
rect 7055 11648 7932 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 8864 11676 8892 11707
rect 9030 11704 9036 11716
rect 9088 11744 9094 11756
rect 9088 11716 9674 11744
rect 9088 11704 9094 11716
rect 8536 11648 8892 11676
rect 8536 11636 8542 11648
rect 8938 11636 8944 11688
rect 8996 11636 9002 11688
rect 9646 11676 9674 11716
rect 9858 11704 9864 11756
rect 9916 11704 9922 11756
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 9968 11676 9996 11707
rect 10042 11704 10048 11756
rect 10100 11704 10106 11756
rect 10226 11704 10232 11756
rect 10284 11704 10290 11756
rect 10502 11704 10508 11756
rect 10560 11704 10566 11756
rect 10594 11704 10600 11756
rect 10652 11744 10658 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 10652 11716 10701 11744
rect 10652 11704 10658 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 9646 11648 9996 11676
rect 10134 11636 10140 11688
rect 10192 11676 10198 11688
rect 10888 11676 10916 11707
rect 11514 11704 11520 11756
rect 11572 11744 11578 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11572 11716 11713 11744
rect 11572 11704 11578 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 12124 11716 12265 11744
rect 12124 11704 12130 11716
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 12526 11704 12532 11756
rect 12584 11704 12590 11756
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11742 12679 11747
rect 12894 11742 12900 11756
rect 12667 11714 12900 11742
rect 12667 11713 12679 11714
rect 12621 11707 12679 11713
rect 12894 11704 12900 11714
rect 12952 11704 12958 11756
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 13648 11753 13676 11852
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 14550 11880 14556 11892
rect 14047 11852 14556 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 14826 11840 14832 11892
rect 14884 11840 14890 11892
rect 16316 11784 16896 11812
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 13044 11716 13093 11744
rect 13044 11704 13050 11716
rect 13081 11713 13093 11716
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11744 13691 11747
rect 14182 11744 14188 11756
rect 13679 11716 14188 11744
rect 13679 11713 13691 11716
rect 13633 11707 13691 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 15194 11744 15200 11756
rect 15059 11716 15200 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 11974 11676 11980 11688
rect 10192 11648 10916 11676
rect 10980 11648 11980 11676
rect 10192 11636 10198 11648
rect 6546 11568 6552 11620
rect 6604 11608 6610 11620
rect 7193 11611 7251 11617
rect 7193 11608 7205 11611
rect 6604 11580 7205 11608
rect 6604 11568 6610 11580
rect 7193 11577 7205 11580
rect 7239 11577 7251 11611
rect 7193 11571 7251 11577
rect 7653 11611 7711 11617
rect 7653 11577 7665 11611
rect 7699 11608 7711 11611
rect 10980 11608 11008 11648
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 12361 11648 13952 11676
rect 7699 11580 11008 11608
rect 11057 11611 11115 11617
rect 7699 11577 7711 11580
rect 7653 11571 7711 11577
rect 11057 11577 11069 11611
rect 11103 11608 11115 11611
rect 12361 11608 12389 11648
rect 13814 11608 13820 11620
rect 11103 11580 12389 11608
rect 12452 11580 13820 11608
rect 11103 11577 11115 11580
rect 11057 11571 11115 11577
rect 2041 11543 2099 11549
rect 2041 11509 2053 11543
rect 2087 11540 2099 11543
rect 2222 11540 2228 11552
rect 2087 11512 2228 11540
rect 2087 11509 2099 11512
rect 2041 11503 2099 11509
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 3326 11500 3332 11552
rect 3384 11500 3390 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4249 11543 4307 11549
rect 4249 11540 4261 11543
rect 4120 11512 4261 11540
rect 4120 11500 4126 11512
rect 4249 11509 4261 11512
rect 4295 11509 4307 11543
rect 4249 11503 4307 11509
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 8168 11512 9597 11540
rect 8168 11500 8174 11512
rect 9585 11509 9597 11512
rect 9631 11540 9643 11543
rect 10594 11540 10600 11552
rect 9631 11512 10600 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 10928 11512 11805 11540
rect 10928 11500 10934 11512
rect 11793 11509 11805 11512
rect 11839 11540 11851 11543
rect 12452 11540 12480 11580
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 13924 11608 13952 11648
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 15028 11676 15056 11707
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 14056 11648 15056 11676
rect 14056 11636 14062 11648
rect 16316 11608 16344 11784
rect 16868 11753 16896 11784
rect 16393 11747 16451 11753
rect 16393 11713 16405 11747
rect 16439 11713 16451 11747
rect 16393 11707 16451 11713
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11744 16911 11747
rect 17218 11744 17224 11756
rect 16899 11716 17224 11744
rect 16899 11713 16911 11716
rect 16853 11707 16911 11713
rect 16408 11676 16436 11707
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17402 11704 17408 11756
rect 17460 11704 17466 11756
rect 17420 11676 17448 11704
rect 16408 11648 17448 11676
rect 13924 11580 16344 11608
rect 11839 11512 12480 11540
rect 13173 11543 13231 11549
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 13538 11540 13544 11552
rect 13219 11512 13544 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 15194 11540 15200 11552
rect 14424 11512 15200 11540
rect 14424 11500 14430 11512
rect 15194 11500 15200 11512
rect 15252 11540 15258 11552
rect 15562 11540 15568 11552
rect 15252 11512 15568 11540
rect 15252 11500 15258 11512
rect 15562 11500 15568 11512
rect 15620 11540 15626 11552
rect 15930 11540 15936 11552
rect 15620 11512 15936 11540
rect 15620 11500 15626 11512
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16206 11500 16212 11552
rect 16264 11500 16270 11552
rect 17405 11543 17463 11549
rect 17405 11509 17417 11543
rect 17451 11540 17463 11543
rect 18138 11540 18144 11552
rect 17451 11512 18144 11540
rect 17451 11509 17463 11512
rect 17405 11503 17463 11509
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 1104 11450 18860 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 18860 11450
rect 1104 11376 18860 11398
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5074 11336 5080 11348
rect 4663 11308 5080 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 6641 11339 6699 11345
rect 6641 11305 6653 11339
rect 6687 11336 6699 11339
rect 6730 11336 6736 11348
rect 6687 11308 6736 11336
rect 6687 11305 6699 11308
rect 6641 11299 6699 11305
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 8113 11339 8171 11345
rect 8113 11305 8125 11339
rect 8159 11336 8171 11339
rect 8754 11336 8760 11348
rect 8159 11308 8760 11336
rect 8159 11305 8171 11308
rect 8113 11299 8171 11305
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 8956 11308 10609 11336
rect 4706 11228 4712 11280
rect 4764 11268 4770 11280
rect 8956 11268 8984 11308
rect 10597 11305 10609 11308
rect 10643 11336 10655 11339
rect 10643 11308 11652 11336
rect 10643 11305 10655 11308
rect 10597 11299 10655 11305
rect 4764 11240 8984 11268
rect 9033 11271 9091 11277
rect 4764 11228 4770 11240
rect 9033 11237 9045 11271
rect 9079 11268 9091 11271
rect 10137 11271 10195 11277
rect 10137 11268 10149 11271
rect 9079 11240 10149 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 10137 11237 10149 11240
rect 10183 11268 10195 11271
rect 11624 11268 11652 11308
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 12618 11336 12624 11348
rect 11756 11308 12624 11336
rect 11756 11296 11762 11308
rect 12618 11296 12624 11308
rect 12676 11336 12682 11348
rect 13170 11336 13176 11348
rect 12676 11308 13176 11336
rect 12676 11296 12682 11308
rect 13170 11296 13176 11308
rect 13228 11336 13234 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13228 11308 13277 11336
rect 13228 11296 13234 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 17310 11336 17316 11348
rect 13412 11308 15608 11336
rect 13412 11296 13418 11308
rect 15470 11268 15476 11280
rect 10183 11240 11560 11268
rect 11624 11240 15476 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 1765 11203 1823 11209
rect 1765 11200 1777 11203
rect 1544 11172 1777 11200
rect 1544 11160 1550 11172
rect 1765 11169 1777 11172
rect 1811 11169 1823 11203
rect 1765 11163 1823 11169
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7742 11200 7748 11212
rect 7055 11172 7748 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 8570 11160 8576 11212
rect 8628 11160 8634 11212
rect 8665 11203 8723 11209
rect 8665 11169 8677 11203
rect 8711 11200 8723 11203
rect 9122 11200 9128 11212
rect 8711 11172 9128 11200
rect 8711 11169 8723 11172
rect 8665 11163 8723 11169
rect 9122 11160 9128 11172
rect 9180 11200 9186 11212
rect 9306 11200 9312 11212
rect 9180 11172 9312 11200
rect 9180 11160 9186 11172
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11200 9551 11203
rect 9582 11200 9588 11212
rect 9539 11172 9588 11200
rect 9539 11169 9551 11172
rect 9493 11163 9551 11169
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 10686 11200 10692 11212
rect 9692 11172 10692 11200
rect 2958 11092 2964 11144
rect 3016 11092 3022 11144
rect 3510 11092 3516 11144
rect 3568 11092 3574 11144
rect 4062 11092 4068 11144
rect 4120 11092 4126 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 5810 11132 5816 11144
rect 4663 11104 5816 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 5972 11135 6030 11141
rect 5972 11101 5984 11135
rect 6018 11132 6030 11135
rect 6546 11132 6552 11144
rect 6018 11104 6552 11132
rect 6018 11101 6030 11104
rect 5972 11095 6030 11101
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 6822 11092 6828 11144
rect 6880 11092 6886 11144
rect 7098 11092 7104 11144
rect 7156 11092 7162 11144
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 8076 11104 8125 11132
rect 8076 11092 8082 11104
rect 8113 11101 8125 11104
rect 8159 11101 8171 11135
rect 8369 11135 8427 11141
rect 8369 11132 8381 11135
rect 8113 11095 8171 11101
rect 8358 11101 8381 11132
rect 8415 11101 8427 11135
rect 8358 11095 8427 11101
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 2222 11024 2228 11076
rect 2280 11024 2286 11076
rect 2314 11024 2320 11076
rect 2372 11024 2378 11076
rect 3418 11024 3424 11076
rect 3476 11024 3482 11076
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 8358 11064 8386 11095
rect 7064 11036 8386 11064
rect 9048 11064 9076 11095
rect 9214 11092 9220 11144
rect 9272 11092 9278 11144
rect 9490 11064 9496 11076
rect 9048 11036 9496 11064
rect 7064 11024 7070 11036
rect 9490 11024 9496 11036
rect 9548 11024 9554 11076
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 6043 10999 6101 11005
rect 6043 10996 6055 10999
rect 5592 10968 6055 10996
rect 5592 10956 5598 10968
rect 6043 10965 6055 10968
rect 6089 10965 6101 10999
rect 6043 10959 6101 10965
rect 8478 10956 8484 11008
rect 8536 10956 8542 11008
rect 8938 10956 8944 11008
rect 8996 10996 9002 11008
rect 9692 10996 9720 11172
rect 10686 11160 10692 11172
rect 10744 11200 10750 11212
rect 11532 11209 11560 11240
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 15580 11268 15608 11308
rect 16132 11308 17316 11336
rect 16022 11268 16028 11280
rect 15580 11240 16028 11268
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 11517 11203 11575 11209
rect 10744 11172 10916 11200
rect 10744 11160 10750 11172
rect 9766 11092 9772 11144
rect 9824 11092 9830 11144
rect 9950 11092 9956 11144
rect 10008 11092 10014 11144
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11132 10287 11135
rect 10410 11132 10416 11144
rect 10275 11104 10416 11132
rect 10275 11101 10287 11104
rect 10229 11095 10287 11101
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 10888 11141 10916 11172
rect 11517 11169 11529 11203
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 13136 11172 14565 11200
rect 13136 11160 13142 11172
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 15286 11200 15292 11212
rect 14553 11163 14611 11169
rect 14936 11172 15292 11200
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11296 11104 11713 11132
rect 11296 11092 11302 11104
rect 11701 11101 11713 11104
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11848 11104 11897 11132
rect 11848 11092 11854 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 12250 11092 12256 11144
rect 12308 11092 12314 11144
rect 12346 11135 12404 11141
rect 12346 11101 12358 11135
rect 12392 11126 12404 11135
rect 12434 11126 12440 11144
rect 12392 11101 12440 11126
rect 12346 11098 12440 11101
rect 12346 11095 12404 11098
rect 12434 11092 12440 11098
rect 12492 11092 12498 11144
rect 14734 11092 14740 11144
rect 14792 11092 14798 11144
rect 14936 11141 14964 11172
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 16132 11200 16160 11308
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 18141 11271 18199 11277
rect 18141 11268 18153 11271
rect 16264 11240 18153 11268
rect 16264 11228 16270 11240
rect 18141 11237 18153 11240
rect 18187 11237 18199 11271
rect 18141 11231 18199 11237
rect 17773 11203 17831 11209
rect 17773 11200 17785 11203
rect 15611 11172 16160 11200
rect 16408 11172 17785 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 15194 11092 15200 11144
rect 15252 11092 15258 11144
rect 15746 11092 15752 11144
rect 15804 11092 15810 11144
rect 16025 11135 16083 11141
rect 16025 11101 16037 11135
rect 16071 11132 16083 11135
rect 16298 11132 16304 11144
rect 16071 11104 16304 11132
rect 16071 11101 16083 11104
rect 16025 11095 16083 11101
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 16408 11141 16436 11172
rect 17773 11169 17785 11172
rect 17819 11169 17831 11203
rect 17773 11163 17831 11169
rect 16393 11135 16451 11141
rect 16393 11101 16405 11135
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11132 17003 11135
rect 17402 11132 17408 11144
rect 16991 11104 17408 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 9861 11067 9919 11073
rect 9861 11033 9873 11067
rect 9907 11064 9919 11067
rect 11606 11064 11612 11076
rect 9907 11036 11612 11064
rect 9907 11033 9919 11036
rect 9861 11027 9919 11033
rect 11606 11024 11612 11036
rect 11664 11024 11670 11076
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 12636 11036 13093 11064
rect 8996 10968 9720 10996
rect 8996 10956 9002 10968
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 11330 10996 11336 11008
rect 11112 10968 11336 10996
rect 11112 10956 11118 10968
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 11790 10956 11796 11008
rect 11848 10996 11854 11008
rect 12636 10996 12664 11036
rect 13081 11033 13093 11036
rect 13127 11033 13139 11067
rect 13630 11064 13636 11076
rect 13081 11027 13139 11033
rect 13188 11036 13636 11064
rect 11848 10968 12664 10996
rect 11848 10956 11854 10968
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13188 10996 13216 11036
rect 12952 10968 13216 10996
rect 12952 10956 12958 10968
rect 13262 10956 13268 11008
rect 13320 11005 13326 11008
rect 13464 11005 13492 11036
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 14829 11067 14887 11073
rect 14829 11033 14841 11067
rect 14875 11033 14887 11067
rect 14829 11027 14887 11033
rect 15059 11067 15117 11073
rect 15059 11033 15071 11067
rect 15105 11064 15117 11067
rect 15838 11064 15844 11076
rect 15105 11036 15844 11064
rect 15105 11033 15117 11036
rect 15059 11027 15117 11033
rect 13320 10999 13339 11005
rect 13327 10965 13339 10999
rect 13320 10959 13339 10965
rect 13449 10999 13507 11005
rect 13449 10965 13461 10999
rect 13495 10965 13507 10999
rect 14844 10996 14872 11027
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 16114 11024 16120 11076
rect 16172 11064 16178 11076
rect 16408 11064 16436 11095
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 16172 11036 16436 11064
rect 16853 11067 16911 11073
rect 16172 11024 16178 11036
rect 16853 11033 16865 11067
rect 16899 11064 16911 11067
rect 18046 11064 18052 11076
rect 16899 11036 18052 11064
rect 16899 11033 16911 11036
rect 16853 11027 16911 11033
rect 18046 11024 18052 11036
rect 18104 11064 18110 11076
rect 18104 11036 18184 11064
rect 18104 11024 18110 11036
rect 15194 10996 15200 11008
rect 14844 10968 15200 10996
rect 13449 10959 13507 10965
rect 13320 10956 13326 10959
rect 15194 10956 15200 10968
rect 15252 10996 15258 11008
rect 15654 10996 15660 11008
rect 15252 10968 15660 10996
rect 15252 10956 15258 10968
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 15930 10956 15936 11008
rect 15988 10956 15994 11008
rect 18156 11005 18184 11036
rect 18141 10999 18199 11005
rect 18141 10965 18153 10999
rect 18187 10965 18199 10999
rect 18141 10959 18199 10965
rect 1104 10906 18860 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 16214 10906
rect 16266 10854 16278 10906
rect 16330 10854 16342 10906
rect 16394 10854 16406 10906
rect 16458 10854 16470 10906
rect 16522 10854 18860 10906
rect 1104 10832 18860 10854
rect 2314 10752 2320 10804
rect 2372 10801 2378 10804
rect 2372 10795 2421 10801
rect 2372 10761 2375 10795
rect 2409 10761 2421 10795
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 2372 10755 2421 10761
rect 2746 10764 3249 10792
rect 2372 10752 2378 10755
rect 2292 10659 2350 10665
rect 2292 10625 2304 10659
rect 2338 10656 2350 10659
rect 2746 10656 2774 10764
rect 3237 10761 3249 10764
rect 3283 10792 3295 10795
rect 3418 10792 3424 10804
rect 3283 10764 3424 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 8110 10792 8116 10804
rect 3936 10764 8116 10792
rect 3936 10752 3942 10764
rect 4985 10727 5043 10733
rect 4985 10693 4997 10727
rect 5031 10724 5043 10727
rect 5534 10724 5540 10736
rect 5031 10696 5540 10724
rect 5031 10693 5043 10696
rect 4985 10687 5043 10693
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 6748 10733 6776 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8665 10795 8723 10801
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 9766 10792 9772 10804
rect 8711 10764 9772 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10008 10764 10149 10792
rect 10008 10752 10014 10764
rect 10137 10761 10149 10764
rect 10183 10792 10195 10795
rect 10226 10792 10232 10804
rect 10183 10764 10232 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 10413 10795 10471 10801
rect 10413 10761 10425 10795
rect 10459 10792 10471 10795
rect 10502 10792 10508 10804
rect 10459 10764 10508 10792
rect 10459 10761 10471 10764
rect 10413 10755 10471 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 10594 10752 10600 10804
rect 10652 10792 10658 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 10652 10764 11897 10792
rect 10652 10752 10658 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12802 10792 12808 10804
rect 12032 10764 12808 10792
rect 12032 10752 12038 10764
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13909 10795 13967 10801
rect 13909 10761 13921 10795
rect 13955 10792 13967 10795
rect 14734 10792 14740 10804
rect 13955 10764 14740 10792
rect 13955 10761 13967 10764
rect 13909 10755 13967 10761
rect 14734 10752 14740 10764
rect 14792 10792 14798 10804
rect 14792 10764 15148 10792
rect 14792 10752 14798 10764
rect 6733 10727 6791 10733
rect 6733 10693 6745 10727
rect 6779 10693 6791 10727
rect 9858 10724 9864 10736
rect 6733 10687 6791 10693
rect 8956 10696 9864 10724
rect 2338 10628 2774 10656
rect 3237 10659 3295 10665
rect 2338 10625 2350 10628
rect 2292 10619 2350 10625
rect 3237 10625 3249 10659
rect 3283 10656 3295 10659
rect 3326 10656 3332 10668
rect 3283 10628 3332 10656
rect 3283 10625 3295 10628
rect 3237 10619 3295 10625
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4212 10628 4445 10656
rect 4212 10616 4218 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10656 4951 10659
rect 5074 10656 5080 10668
rect 4939 10628 5080 10656
rect 4939 10625 4951 10628
rect 4893 10619 4951 10625
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5328 10659 5386 10665
rect 5328 10625 5340 10659
rect 5374 10656 5386 10659
rect 5902 10656 5908 10668
rect 5374 10628 5908 10656
rect 5374 10625 5386 10628
rect 5328 10619 5386 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 2869 10591 2927 10597
rect 2869 10557 2881 10591
rect 2915 10588 2927 10591
rect 2958 10588 2964 10600
rect 2915 10560 2964 10588
rect 2915 10557 2927 10560
rect 2869 10551 2927 10557
rect 2958 10548 2964 10560
rect 3016 10588 3022 10600
rect 4798 10588 4804 10600
rect 3016 10560 4804 10588
rect 3016 10548 3022 10560
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 6564 10588 6592 10619
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 6825 10659 6883 10665
rect 6696 10655 6776 10656
rect 6825 10655 6837 10659
rect 6696 10628 6837 10655
rect 6696 10616 6702 10628
rect 6748 10627 6837 10628
rect 6825 10625 6837 10627
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 7650 10665 7656 10668
rect 7621 10659 7656 10665
rect 7621 10625 7633 10659
rect 7621 10619 7656 10625
rect 7650 10616 7656 10619
rect 7708 10616 7714 10668
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 8110 10656 8116 10668
rect 7800 10628 8116 10656
rect 7800 10616 7806 10628
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 8956 10665 8984 10696
rect 9858 10684 9864 10696
rect 9916 10684 9922 10736
rect 11330 10724 11336 10736
rect 10612 10696 11336 10724
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 9950 10656 9956 10668
rect 9548 10628 9956 10656
rect 9548 10616 9554 10628
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 10502 10656 10508 10668
rect 10183 10628 10508 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10612 10665 10640 10696
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 14826 10724 14832 10736
rect 11808 10696 14832 10724
rect 10598 10659 10656 10665
rect 10598 10625 10610 10659
rect 10644 10625 10656 10659
rect 10598 10619 10656 10625
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10656 10747 10659
rect 10965 10659 11023 10665
rect 10735 10628 10824 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 7466 10588 7472 10600
rect 6564 10560 7472 10588
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 8846 10588 8852 10600
rect 7883 10560 8852 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9048 10588 9076 10616
rect 10612 10588 10640 10619
rect 10796 10588 10824 10628
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11606 10656 11612 10668
rect 11011 10628 11612 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 9048 10560 10640 10588
rect 10704 10560 10824 10588
rect 3970 10480 3976 10532
rect 4028 10520 4034 10532
rect 10134 10520 10140 10532
rect 4028 10492 10140 10520
rect 4028 10480 4034 10492
rect 10134 10480 10140 10492
rect 10192 10480 10198 10532
rect 10410 10480 10416 10532
rect 10468 10520 10474 10532
rect 10704 10520 10732 10560
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 11808 10520 11836 10696
rect 14826 10684 14832 10696
rect 14884 10684 14890 10736
rect 15120 10733 15148 10764
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 15712 10764 16221 10792
rect 15712 10752 15718 10764
rect 16209 10761 16221 10764
rect 16255 10761 16267 10795
rect 16209 10755 16267 10761
rect 17221 10795 17279 10801
rect 17221 10761 17233 10795
rect 17267 10792 17279 10795
rect 17954 10792 17960 10804
rect 17267 10764 17960 10792
rect 17267 10761 17279 10764
rect 17221 10755 17279 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 15105 10727 15163 10733
rect 15105 10693 15117 10727
rect 15151 10693 15163 10727
rect 15105 10687 15163 10693
rect 15194 10684 15200 10736
rect 15252 10724 15258 10736
rect 15378 10733 15384 10736
rect 15335 10727 15384 10733
rect 15252 10696 15297 10724
rect 15252 10684 15258 10696
rect 15335 10693 15347 10727
rect 15381 10693 15384 10727
rect 15335 10687 15384 10693
rect 15378 10684 15384 10687
rect 15436 10684 15442 10736
rect 15470 10684 15476 10736
rect 15528 10724 15534 10736
rect 15841 10727 15899 10733
rect 15841 10724 15853 10727
rect 15528 10696 15853 10724
rect 15528 10684 15534 10696
rect 15841 10693 15853 10696
rect 15887 10693 15899 10727
rect 15841 10687 15899 10693
rect 16071 10693 16129 10699
rect 16071 10690 16083 10693
rect 12066 10616 12072 10668
rect 12124 10616 12130 10668
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10625 12311 10659
rect 12253 10619 12311 10625
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12713 10659 12771 10665
rect 12713 10625 12725 10659
rect 12759 10656 12771 10659
rect 12802 10656 12808 10668
rect 12759 10628 12808 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 12268 10588 12296 10619
rect 11940 10560 12296 10588
rect 11940 10548 11946 10560
rect 10468 10492 10732 10520
rect 11072 10492 11836 10520
rect 12360 10520 12388 10619
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 13170 10616 13176 10668
rect 13228 10616 13234 10668
rect 13354 10616 13360 10668
rect 13412 10616 13418 10668
rect 13538 10616 13544 10668
rect 13596 10616 13602 10668
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 13906 10656 13912 10668
rect 13771 10628 13912 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14274 10656 14280 10668
rect 14231 10628 14280 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 15010 10616 15016 10668
rect 15068 10616 15074 10668
rect 16056 10659 16083 10690
rect 16117 10659 16129 10693
rect 18138 10684 18144 10736
rect 18196 10684 18202 10736
rect 18230 10684 18236 10736
rect 18288 10684 18294 10736
rect 16056 10656 16129 10659
rect 15120 10653 16129 10656
rect 15120 10628 16084 10653
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 13449 10591 13507 10597
rect 13449 10588 13461 10591
rect 12584 10560 13461 10588
rect 12584 10548 12590 10560
rect 13449 10557 13461 10560
rect 13495 10588 13507 10591
rect 13630 10588 13636 10600
rect 13495 10560 13636 10588
rect 13495 10557 13507 10560
rect 13449 10551 13507 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15120 10588 15148 10628
rect 17218 10616 17224 10668
rect 17276 10656 17282 10668
rect 17681 10659 17739 10665
rect 17681 10656 17693 10659
rect 17276 10628 17693 10656
rect 17276 10616 17282 10628
rect 17681 10625 17693 10628
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 14976 10560 15148 10588
rect 14976 10548 14982 10560
rect 15194 10548 15200 10600
rect 15252 10588 15258 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 15252 10560 15485 10588
rect 15252 10548 15258 10560
rect 15473 10557 15485 10560
rect 15519 10588 15531 10591
rect 15930 10588 15936 10600
rect 15519 10560 15936 10588
rect 15519 10557 15531 10560
rect 15473 10551 15531 10557
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16758 10548 16764 10600
rect 16816 10588 16822 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16816 10560 16865 10588
rect 16816 10548 16822 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 16853 10551 16911 10557
rect 12618 10520 12624 10532
rect 12360 10492 12624 10520
rect 10468 10480 10474 10492
rect 4706 10412 4712 10464
rect 4764 10452 4770 10464
rect 5399 10455 5457 10461
rect 5399 10452 5411 10455
rect 4764 10424 5411 10452
rect 4764 10412 4770 10424
rect 5399 10421 5411 10424
rect 5445 10421 5457 10455
rect 5399 10415 5457 10421
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 7101 10455 7159 10461
rect 7101 10452 7113 10455
rect 5592 10424 7113 10452
rect 5592 10412 5598 10424
rect 7101 10421 7113 10424
rect 7147 10421 7159 10455
rect 7101 10415 7159 10421
rect 7374 10412 7380 10464
rect 7432 10412 7438 10464
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 11072 10452 11100 10492
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 13078 10480 13084 10532
rect 13136 10520 13142 10532
rect 13262 10520 13268 10532
rect 13136 10492 13268 10520
rect 13136 10480 13142 10492
rect 13262 10480 13268 10492
rect 13320 10520 13326 10532
rect 14829 10523 14887 10529
rect 13320 10492 14412 10520
rect 13320 10480 13326 10492
rect 8444 10424 11100 10452
rect 8444 10412 8450 10424
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 12250 10452 12256 10464
rect 11204 10424 12256 10452
rect 11204 10412 11210 10424
rect 12250 10412 12256 10424
rect 12308 10452 12314 10464
rect 12710 10452 12716 10464
rect 12308 10424 12716 10452
rect 12308 10412 12314 10424
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 13780 10424 14289 10452
rect 13780 10412 13786 10424
rect 14277 10421 14289 10424
rect 14323 10421 14335 10455
rect 14384 10452 14412 10492
rect 14829 10489 14841 10523
rect 14875 10520 14887 10523
rect 16114 10520 16120 10532
rect 14875 10492 16120 10520
rect 14875 10489 14887 10492
rect 14829 10483 14887 10489
rect 16114 10480 16120 10492
rect 16172 10480 16178 10532
rect 17218 10480 17224 10532
rect 17276 10480 17282 10532
rect 16025 10455 16083 10461
rect 16025 10452 16037 10455
rect 14384 10424 16037 10452
rect 14277 10415 14335 10421
rect 16025 10421 16037 10424
rect 16071 10421 16083 10455
rect 16025 10415 16083 10421
rect 1104 10362 18860 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 18860 10362
rect 1104 10288 18860 10310
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10248 4583 10251
rect 8938 10248 8944 10260
rect 4571 10220 8248 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 5261 10183 5319 10189
rect 5261 10149 5273 10183
rect 5307 10180 5319 10183
rect 5721 10183 5779 10189
rect 5721 10180 5733 10183
rect 5307 10152 5733 10180
rect 5307 10149 5319 10152
rect 5261 10143 5319 10149
rect 5721 10149 5733 10152
rect 5767 10149 5779 10183
rect 5721 10143 5779 10149
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 7745 10183 7803 10189
rect 7745 10180 7757 10183
rect 7708 10152 7757 10180
rect 7708 10140 7714 10152
rect 7745 10149 7757 10152
rect 7791 10149 7803 10183
rect 7745 10143 7803 10149
rect 7926 10140 7932 10192
rect 7984 10140 7990 10192
rect 7374 10112 7380 10124
rect 6380 10084 7380 10112
rect 2222 10004 2228 10056
rect 2280 10044 2286 10056
rect 2352 10047 2410 10053
rect 2352 10044 2364 10047
rect 2280 10016 2364 10044
rect 2280 10004 2286 10016
rect 2352 10013 2364 10016
rect 2398 10013 2410 10047
rect 2352 10007 2410 10013
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5534 10044 5540 10056
rect 4939 10016 5540 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 6380 10053 6408 10084
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 8220 10112 8248 10220
rect 8404 10220 8944 10248
rect 8404 10189 8432 10220
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9306 10248 9312 10260
rect 9079 10220 9312 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9490 10208 9496 10260
rect 9548 10208 9554 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10226 10248 10232 10260
rect 10183 10220 10232 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 10520 10220 10916 10248
rect 8389 10183 8447 10189
rect 8389 10149 8401 10183
rect 8435 10149 8447 10183
rect 9766 10180 9772 10192
rect 8389 10143 8447 10149
rect 8588 10152 9772 10180
rect 8588 10112 8616 10152
rect 9766 10140 9772 10152
rect 9824 10140 9830 10192
rect 10410 10140 10416 10192
rect 10468 10140 10474 10192
rect 8220 10084 8616 10112
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 10428 10112 10456 10140
rect 9088 10084 9536 10112
rect 9088 10072 9094 10084
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5868 10016 5917 10044
rect 5868 10004 5874 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 8018 10044 8024 10056
rect 6687 10016 8024 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 8386 10004 8392 10056
rect 8444 10004 8450 10056
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 8662 10044 8668 10056
rect 8619 10016 8668 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 9214 10004 9220 10056
rect 9272 10004 9278 10056
rect 9369 10047 9427 10053
rect 9369 10013 9381 10047
rect 9415 10044 9427 10047
rect 9415 10040 9444 10044
rect 9508 10040 9536 10084
rect 10244 10084 10456 10112
rect 9415 10013 9536 10040
rect 9369 10012 9536 10013
rect 9369 10007 9427 10012
rect 9582 10004 9588 10056
rect 9640 10004 9646 10056
rect 10134 10004 10140 10056
rect 10192 10004 10198 10056
rect 4433 9979 4491 9985
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 4614 9976 4620 9988
rect 4479 9948 4620 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 4798 9936 4804 9988
rect 4856 9976 4862 9988
rect 7469 9979 7527 9985
rect 4856 9948 7328 9976
rect 4856 9936 4862 9948
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 2455 9911 2513 9917
rect 2455 9908 2467 9911
rect 2096 9880 2467 9908
rect 2096 9868 2102 9880
rect 2455 9877 2467 9880
rect 2501 9877 2513 9911
rect 2455 9871 2513 9877
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 5902 9908 5908 9920
rect 5307 9880 5908 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 6178 9868 6184 9920
rect 6236 9868 6242 9920
rect 6549 9911 6607 9917
rect 6549 9877 6561 9911
rect 6595 9908 6607 9911
rect 7190 9908 7196 9920
rect 6595 9880 7196 9908
rect 6595 9877 6607 9880
rect 6549 9871 6607 9877
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7300 9908 7328 9948
rect 7469 9945 7481 9979
rect 7515 9976 7527 9979
rect 7558 9976 7564 9988
rect 7515 9948 7564 9976
rect 7515 9945 7527 9948
rect 7469 9939 7527 9945
rect 7558 9936 7564 9948
rect 7616 9936 7622 9988
rect 9766 9976 9772 9988
rect 9508 9948 9772 9976
rect 8754 9908 8760 9920
rect 7300 9880 8760 9908
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 9508 9908 9536 9948
rect 9766 9936 9772 9948
rect 9824 9976 9830 9988
rect 10244 9976 10272 10084
rect 10315 10047 10373 10053
rect 10315 10013 10327 10047
rect 10361 10044 10373 10047
rect 10520 10044 10548 10220
rect 10888 10180 10916 10220
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 11940 10220 12173 10248
rect 11940 10208 11946 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 12618 10208 12624 10260
rect 12676 10208 12682 10260
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 12768 10220 13553 10248
rect 12768 10208 12774 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 13541 10211 13599 10217
rect 15286 10208 15292 10260
rect 15344 10208 15350 10260
rect 11422 10180 11428 10192
rect 10888 10152 11428 10180
rect 11422 10140 11428 10152
rect 11480 10140 11486 10192
rect 12636 10180 12664 10208
rect 12636 10152 12940 10180
rect 12618 10112 12624 10124
rect 10796 10084 12624 10112
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10361 10016 10456 10044
rect 10520 10016 10609 10044
rect 10361 10013 10373 10016
rect 10315 10007 10373 10013
rect 10428 9988 10456 10016
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 10796 10053 10824 10084
rect 10781 10047 10839 10053
rect 10781 10044 10793 10047
rect 10744 10016 10793 10044
rect 10744 10004 10750 10016
rect 10781 10013 10793 10016
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 11624 10053 11652 10084
rect 12618 10072 12624 10084
rect 12676 10112 12682 10124
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12676 10084 12817 10112
rect 12676 10072 12682 10084
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 12912 10112 12940 10152
rect 13078 10140 13084 10192
rect 13136 10140 13142 10192
rect 13188 10152 14596 10180
rect 13188 10112 13216 10152
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 12912 10084 13216 10112
rect 13372 10084 14473 10112
rect 12805 10075 12863 10081
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 11790 10004 11796 10056
rect 11848 10044 11854 10056
rect 12069 10047 12127 10053
rect 12069 10044 12081 10047
rect 11848 10016 12081 10044
rect 11848 10004 11854 10016
rect 12069 10013 12081 10016
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13170 10044 13176 10056
rect 12952 10016 13176 10044
rect 12952 10004 12958 10016
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 13372 10053 13400 10084
rect 14461 10081 14473 10084
rect 14507 10081 14519 10115
rect 14568 10112 14596 10152
rect 15010 10140 15016 10192
rect 15068 10180 15074 10192
rect 15657 10183 15715 10189
rect 15657 10180 15669 10183
rect 15068 10152 15669 10180
rect 15068 10140 15074 10152
rect 15657 10149 15669 10152
rect 15703 10149 15715 10183
rect 15657 10143 15715 10149
rect 17129 10183 17187 10189
rect 17129 10149 17141 10183
rect 17175 10180 17187 10183
rect 17954 10180 17960 10192
rect 17175 10152 17960 10180
rect 17175 10149 17187 10152
rect 17129 10143 17187 10149
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 17034 10112 17040 10124
rect 14568 10084 17040 10112
rect 14461 10075 14519 10081
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10044 13691 10047
rect 13814 10044 13820 10056
rect 13679 10016 13820 10044
rect 13679 10013 13691 10016
rect 13633 10007 13691 10013
rect 9824 9948 10272 9976
rect 9824 9936 9830 9948
rect 10410 9936 10416 9988
rect 10468 9936 10474 9988
rect 10502 9936 10508 9988
rect 10560 9976 10566 9988
rect 12621 9979 12679 9985
rect 10560 9948 10732 9976
rect 10560 9936 10566 9948
rect 9456 9880 9536 9908
rect 9456 9868 9462 9880
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 10594 9908 10600 9920
rect 9640 9880 10600 9908
rect 9640 9868 9646 9880
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 10704 9917 10732 9948
rect 12621 9945 12633 9979
rect 12667 9976 12679 9979
rect 12802 9976 12808 9988
rect 12667 9948 12808 9976
rect 12667 9945 12679 9948
rect 12621 9939 12679 9945
rect 12802 9936 12808 9948
rect 12860 9936 12866 9988
rect 13372 9976 13400 10007
rect 13814 10004 13820 10016
rect 13872 10044 13878 10056
rect 15197 10047 15255 10053
rect 15197 10044 15209 10047
rect 13872 10016 15209 10044
rect 13872 10004 13878 10016
rect 15197 10013 15209 10016
rect 15243 10013 15255 10047
rect 15197 10007 15255 10013
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10044 15347 10047
rect 15654 10044 15660 10056
rect 15335 10016 15660 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 15654 10004 15660 10016
rect 15712 10044 15718 10056
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 15712 10016 15853 10044
rect 15712 10004 15718 10016
rect 15841 10013 15853 10016
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 16758 10004 16764 10056
rect 16816 10004 16822 10056
rect 18049 10047 18107 10053
rect 18049 10013 18061 10047
rect 18095 10044 18107 10047
rect 18138 10044 18144 10056
rect 18095 10016 18144 10044
rect 18095 10013 18107 10016
rect 18049 10007 18107 10013
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 12912 9948 13400 9976
rect 10689 9911 10747 9917
rect 10689 9877 10701 9911
rect 10735 9908 10747 9911
rect 10870 9908 10876 9920
rect 10735 9880 10876 9908
rect 10735 9877 10747 9880
rect 10689 9871 10747 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11514 9868 11520 9920
rect 11572 9868 11578 9920
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 12912 9908 12940 9948
rect 14090 9936 14096 9988
rect 14148 9976 14154 9988
rect 14277 9979 14335 9985
rect 14277 9976 14289 9979
rect 14148 9948 14289 9976
rect 14148 9936 14154 9948
rect 14277 9945 14289 9948
rect 14323 9945 14335 9979
rect 14277 9939 14335 9945
rect 14826 9936 14832 9988
rect 14884 9976 14890 9988
rect 15013 9979 15071 9985
rect 15013 9976 15025 9979
rect 14884 9948 15025 9976
rect 14884 9936 14890 9948
rect 15013 9945 15025 9948
rect 15059 9976 15071 9979
rect 15565 9979 15623 9985
rect 15565 9976 15577 9979
rect 15059 9948 15577 9976
rect 15059 9945 15071 9948
rect 15013 9939 15071 9945
rect 15565 9945 15577 9948
rect 15611 9945 15623 9979
rect 15565 9939 15623 9945
rect 15749 9979 15807 9985
rect 15749 9945 15761 9979
rect 15795 9945 15807 9979
rect 15749 9939 15807 9945
rect 17129 9979 17187 9985
rect 17129 9945 17141 9979
rect 17175 9976 17187 9979
rect 17402 9976 17408 9988
rect 17175 9948 17408 9976
rect 17175 9945 17187 9948
rect 17129 9939 17187 9945
rect 11664 9880 12940 9908
rect 11664 9868 11670 9880
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13906 9908 13912 9920
rect 13136 9880 13912 9908
rect 13136 9868 13142 9880
rect 13906 9868 13912 9880
rect 13964 9908 13970 9920
rect 15764 9908 15792 9939
rect 17402 9936 17408 9948
rect 17460 9976 17466 9988
rect 18233 9979 18291 9985
rect 18233 9976 18245 9979
rect 17460 9948 18245 9976
rect 17460 9936 17466 9948
rect 18233 9945 18245 9948
rect 18279 9945 18291 9979
rect 18233 9939 18291 9945
rect 13964 9880 15792 9908
rect 13964 9868 13970 9880
rect 1104 9818 18860 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 16214 9818
rect 16266 9766 16278 9818
rect 16330 9766 16342 9818
rect 16394 9766 16406 9818
rect 16458 9766 16470 9818
rect 16522 9766 18860 9818
rect 1104 9744 18860 9766
rect 5902 9664 5908 9716
rect 5960 9664 5966 9716
rect 7466 9664 7472 9716
rect 7524 9664 7530 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7616 9676 8248 9704
rect 7616 9664 7622 9676
rect 7285 9639 7343 9645
rect 7285 9605 7297 9639
rect 7331 9636 7343 9639
rect 8021 9639 8079 9645
rect 8021 9636 8033 9639
rect 7331 9608 8033 9636
rect 7331 9605 7343 9608
rect 7285 9599 7343 9605
rect 8021 9605 8033 9608
rect 8067 9605 8079 9639
rect 8220 9636 8248 9676
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 9398 9704 9404 9716
rect 8720 9676 9404 9704
rect 8720 9664 8726 9676
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 11057 9707 11115 9713
rect 11057 9704 11069 9707
rect 10008 9676 11069 9704
rect 10008 9664 10014 9676
rect 11057 9673 11069 9676
rect 11103 9673 11115 9707
rect 11057 9667 11115 9673
rect 12066 9664 12072 9716
rect 12124 9704 12130 9716
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 12124 9676 12173 9704
rect 12124 9664 12130 9676
rect 12161 9673 12173 9676
rect 12207 9673 12219 9707
rect 12894 9704 12900 9716
rect 12161 9667 12219 9673
rect 12406 9676 12900 9704
rect 9214 9636 9220 9648
rect 8220 9608 9220 9636
rect 8021 9599 8079 9605
rect 9214 9596 9220 9608
rect 9272 9636 9278 9648
rect 10686 9636 10692 9648
rect 9272 9608 9352 9636
rect 9272 9596 9278 9608
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 2222 9568 2228 9580
rect 1903 9540 2228 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3145 9571 3203 9577
rect 3145 9568 3157 9571
rect 3108 9540 3157 9568
rect 3108 9528 3114 9540
rect 3145 9537 3157 9540
rect 3191 9537 3203 9571
rect 3145 9531 3203 9537
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 4982 9568 4988 9580
rect 3743 9540 4988 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5534 9528 5540 9580
rect 5592 9528 5598 9580
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 9030 9568 9036 9580
rect 7984 9540 9036 9568
rect 7984 9528 7990 9540
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 9324 9577 9352 9608
rect 9416 9608 10692 9636
rect 9416 9580 9444 9608
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 10889 9639 10947 9645
rect 10889 9636 10901 9639
rect 10796 9608 10901 9636
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 5000 9500 5028 9528
rect 5810 9500 5816 9512
rect 2179 9472 4752 9500
rect 5000 9472 5816 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 2148 9432 2176 9463
rect 1912 9404 2176 9432
rect 3697 9435 3755 9441
rect 1912 9392 1918 9404
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 4614 9432 4620 9444
rect 3743 9404 4620 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 4724 9432 4752 9472
rect 5810 9460 5816 9472
rect 5868 9500 5874 9512
rect 5905 9503 5963 9509
rect 5905 9500 5917 9503
rect 5868 9472 5917 9500
rect 5868 9460 5874 9472
rect 5905 9469 5917 9472
rect 5951 9469 5963 9503
rect 5905 9463 5963 9469
rect 6917 9503 6975 9509
rect 6917 9469 6929 9503
rect 6963 9500 6975 9503
rect 7650 9500 7656 9512
rect 6963 9472 7656 9500
rect 6963 9469 6975 9472
rect 6917 9463 6975 9469
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8570 9500 8576 9512
rect 8067 9472 8576 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9140 9500 9168 9531
rect 9398 9528 9404 9580
rect 9456 9528 9462 9580
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9640 9540 9781 9568
rect 9640 9528 9646 9540
rect 9769 9537 9781 9540
rect 9815 9568 9827 9571
rect 10796 9568 10824 9608
rect 10889 9605 10901 9608
rect 10935 9605 10947 9639
rect 12406 9636 12434 9676
rect 12894 9664 12900 9676
rect 12952 9704 12958 9716
rect 13722 9704 13728 9716
rect 12952 9676 13728 9704
rect 12952 9664 12958 9676
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 15286 9704 15292 9716
rect 14608 9676 15292 9704
rect 14608 9664 14614 9676
rect 15286 9664 15292 9676
rect 15344 9704 15350 9716
rect 15381 9707 15439 9713
rect 15381 9704 15393 9707
rect 15344 9676 15393 9704
rect 15344 9664 15350 9676
rect 15381 9673 15393 9676
rect 15427 9673 15439 9707
rect 16209 9707 16267 9713
rect 16209 9704 16221 9707
rect 15381 9667 15439 9673
rect 15764 9676 16221 9704
rect 10889 9599 10947 9605
rect 11900 9608 12434 9636
rect 11698 9568 11704 9580
rect 9815 9540 11704 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 11900 9577 11928 9608
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 13078 9636 13084 9648
rect 12768 9608 13084 9636
rect 12768 9596 12774 9608
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 14090 9636 14096 9648
rect 13556 9608 14096 9636
rect 13556 9580 13584 9608
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 14182 9596 14188 9648
rect 14240 9596 14246 9648
rect 14369 9639 14427 9645
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 14458 9636 14464 9648
rect 14415 9608 14464 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 15470 9636 15476 9648
rect 14660 9608 15476 9636
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 11974 9528 11980 9580
rect 12032 9568 12038 9580
rect 12032 9540 12434 9568
rect 12032 9528 12038 9540
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9140 9472 10057 9500
rect 10045 9469 10057 9472
rect 10091 9500 10103 9503
rect 12066 9500 12072 9512
rect 10091 9472 12072 9500
rect 10091 9469 10103 9472
rect 10045 9463 10103 9469
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12406 9500 12434 9540
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9568 12955 9571
rect 12986 9568 12992 9580
rect 12943 9540 12992 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 13412 9540 13461 9568
rect 13412 9528 13418 9540
rect 13449 9537 13461 9540
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 13538 9528 13544 9580
rect 13596 9528 13602 9580
rect 13630 9528 13636 9580
rect 13688 9528 13694 9580
rect 14200 9568 14228 9596
rect 14660 9577 14688 9608
rect 15470 9596 15476 9608
rect 15528 9636 15534 9648
rect 15764 9636 15792 9676
rect 16209 9673 16221 9676
rect 16255 9673 16267 9707
rect 16209 9667 16267 9673
rect 15528 9608 15792 9636
rect 15841 9639 15899 9645
rect 15528 9596 15534 9608
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 16758 9636 16764 9648
rect 15887 9608 16764 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 16758 9596 16764 9608
rect 16816 9596 16822 9648
rect 14553 9571 14611 9577
rect 14553 9568 14565 9571
rect 14200 9540 14565 9568
rect 14553 9537 14565 9540
rect 14599 9537 14611 9571
rect 14553 9531 14611 9537
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 15102 9568 15108 9580
rect 14967 9540 15108 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 14844 9500 14872 9531
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 15252 9540 15301 9568
rect 15252 9528 15258 9540
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9537 16359 9571
rect 16301 9531 16359 9537
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9568 16911 9571
rect 17126 9568 17132 9580
rect 16899 9540 17132 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 16040 9500 16068 9531
rect 16316 9500 16344 9531
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 12406 9472 16068 9500
rect 16224 9472 16344 9500
rect 6546 9432 6552 9444
rect 4724 9404 6552 9432
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 7558 9392 7564 9444
rect 7616 9432 7622 9444
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 7616 9404 7849 9432
rect 7616 9392 7622 9404
rect 7837 9401 7849 9404
rect 7883 9401 7895 9435
rect 8849 9435 8907 9441
rect 8849 9432 8861 9435
rect 7837 9395 7895 9401
rect 8036 9404 8861 9432
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 6822 9364 6828 9376
rect 3292 9336 6828 9364
rect 3292 9324 3298 9336
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 8036 9364 8064 9404
rect 8849 9401 8861 9404
rect 8895 9401 8907 9435
rect 10134 9432 10140 9444
rect 8849 9395 8907 9401
rect 10060 9404 10140 9432
rect 7331 9336 8064 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 8996 9336 9873 9364
rect 8996 9324 9002 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 9953 9367 10011 9373
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10060 9364 10088 9404
rect 10134 9392 10140 9404
rect 10192 9392 10198 9444
rect 11882 9392 11888 9444
rect 11940 9432 11946 9444
rect 12713 9435 12771 9441
rect 12713 9432 12725 9435
rect 11940 9404 12725 9432
rect 11940 9392 11946 9404
rect 12713 9401 12725 9404
rect 12759 9401 12771 9435
rect 12713 9395 12771 9401
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9432 12863 9435
rect 13354 9432 13360 9444
rect 12851 9404 13360 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 13446 9392 13452 9444
rect 13504 9432 13510 9444
rect 13630 9432 13636 9444
rect 13504 9404 13636 9432
rect 13504 9392 13510 9404
rect 13630 9392 13636 9404
rect 13688 9392 13694 9444
rect 13817 9435 13875 9441
rect 13817 9401 13829 9435
rect 13863 9432 13875 9435
rect 14918 9432 14924 9444
rect 13863 9404 14924 9432
rect 13863 9401 13875 9404
rect 13817 9395 13875 9401
rect 14918 9392 14924 9404
rect 14976 9392 14982 9444
rect 15746 9432 15752 9444
rect 15028 9404 15752 9432
rect 9999 9336 10088 9364
rect 10873 9367 10931 9373
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10873 9333 10885 9367
rect 10919 9364 10931 9367
rect 11606 9364 11612 9376
rect 10919 9336 11612 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 15028 9364 15056 9404
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 15930 9392 15936 9444
rect 15988 9432 15994 9444
rect 16224 9432 16252 9472
rect 15988 9404 16252 9432
rect 15988 9392 15994 9404
rect 12483 9336 15056 9364
rect 17405 9367 17463 9373
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 17405 9333 17417 9367
rect 17451 9364 17463 9367
rect 17586 9364 17592 9376
rect 17451 9336 17592 9364
rect 17451 9333 17463 9336
rect 17405 9327 17463 9333
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 1104 9274 18860 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 18860 9274
rect 1104 9200 18860 9222
rect 3050 9120 3056 9172
rect 3108 9120 3114 9172
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 7190 9120 7196 9172
rect 7248 9160 7254 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 7248 9132 7941 9160
rect 7248 9120 7254 9132
rect 7929 9129 7941 9132
rect 7975 9129 7987 9163
rect 7929 9123 7987 9129
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9398 9160 9404 9172
rect 9171 9132 9404 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 9769 9163 9827 9169
rect 9769 9129 9781 9163
rect 9815 9160 9827 9163
rect 9858 9160 9864 9172
rect 9815 9132 9864 9160
rect 9815 9129 9827 9132
rect 9769 9123 9827 9129
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 11333 9163 11391 9169
rect 11333 9160 11345 9163
rect 10336 9132 11345 9160
rect 3068 9092 3096 9120
rect 4341 9095 4399 9101
rect 3068 9064 3924 9092
rect 1302 8984 1308 9036
rect 1360 9024 1366 9036
rect 3896 9033 3924 9064
rect 4341 9061 4353 9095
rect 4387 9092 4399 9095
rect 4614 9092 4620 9104
rect 4387 9064 4620 9092
rect 4387 9061 4399 9064
rect 4341 9055 4399 9061
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 7208 9064 9536 9092
rect 3881 9027 3939 9033
rect 1360 8996 3556 9024
rect 1360 8984 1366 8996
rect 1210 8916 1216 8968
rect 1268 8956 1274 8968
rect 2041 8959 2099 8965
rect 1268 8928 1992 8956
rect 1268 8916 1274 8928
rect 1854 8848 1860 8900
rect 1912 8848 1918 8900
rect 1964 8888 1992 8928
rect 2041 8925 2053 8959
rect 2087 8956 2099 8959
rect 2130 8956 2136 8968
rect 2087 8928 2136 8956
rect 2087 8925 2099 8928
rect 2041 8919 2099 8925
rect 2130 8916 2136 8928
rect 2188 8956 2194 8968
rect 2314 8956 2320 8968
rect 2188 8928 2320 8956
rect 2188 8916 2194 8928
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 2516 8888 2544 8919
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3528 8965 3556 8996
rect 3881 8993 3893 9027
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4706 9024 4712 9036
rect 4479 8996 4712 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 5512 8959 5570 8965
rect 5512 8925 5524 8959
rect 5558 8956 5570 8959
rect 6086 8956 6092 8968
rect 5558 8928 6092 8956
rect 5558 8925 5570 8928
rect 5512 8919 5570 8925
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 7098 8916 7104 8968
rect 7156 8916 7162 8968
rect 7208 8965 7236 9064
rect 9508 9036 9536 9064
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 10229 9095 10287 9101
rect 10229 9092 10241 9095
rect 9732 9064 10241 9092
rect 9732 9052 9738 9064
rect 10229 9061 10241 9064
rect 10275 9061 10287 9095
rect 10229 9055 10287 9061
rect 7282 8984 7288 9036
rect 7340 8984 7346 9036
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 7984 8996 8524 9024
rect 7984 8984 7990 8996
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8925 7251 8959
rect 7193 8919 7251 8925
rect 1964 8860 2544 8888
rect 4890 8848 4896 8900
rect 4948 8848 4954 8900
rect 6362 8848 6368 8900
rect 6420 8848 6426 8900
rect 6914 8848 6920 8900
rect 6972 8848 6978 8900
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8820 2559 8823
rect 2958 8820 2964 8832
rect 2547 8792 2964 8820
rect 2547 8789 2559 8792
rect 2501 8783 2559 8789
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3418 8780 3424 8832
rect 3476 8780 3482 8832
rect 5534 8780 5540 8832
rect 5592 8829 5598 8832
rect 5592 8823 5641 8829
rect 5592 8789 5595 8823
rect 5629 8789 5641 8823
rect 5592 8783 5641 8789
rect 5592 8780 5598 8783
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7208 8820 7236 8919
rect 7374 8916 7380 8968
rect 7432 8965 7438 8968
rect 8496 8965 8524 8996
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 10336 9024 10364 9132
rect 11333 9129 11345 9132
rect 11379 9129 11391 9163
rect 11333 9123 11391 9129
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 11756 9132 12081 9160
rect 11756 9120 11762 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12069 9123 12127 9129
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13044 9132 15148 9160
rect 13044 9120 13050 9132
rect 13449 9095 13507 9101
rect 13449 9061 13461 9095
rect 13495 9092 13507 9095
rect 13630 9092 13636 9104
rect 13495 9064 13636 9092
rect 13495 9061 13507 9064
rect 13449 9055 13507 9061
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 14458 9092 14464 9104
rect 13740 9064 14464 9092
rect 10870 9024 10876 9036
rect 9548 8996 10364 9024
rect 10428 8996 10876 9024
rect 9548 8984 9554 8996
rect 7432 8959 7447 8965
rect 7435 8925 7447 8959
rect 7432 8919 7447 8925
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8956 8539 8959
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8527 8928 9045 8956
rect 8527 8925 8539 8928
rect 8481 8919 8539 8925
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 9766 8956 9772 8968
rect 9723 8928 9772 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 7432 8916 7438 8919
rect 7834 8848 7840 8900
rect 7892 8848 7898 8900
rect 8312 8888 8340 8919
rect 8754 8888 8760 8900
rect 8312 8860 8760 8888
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 7156 8792 7236 8820
rect 7156 8780 7162 8792
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 7708 8792 8401 8820
rect 7708 8780 7714 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 9048 8820 9076 8919
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 9950 8956 9956 8968
rect 9907 8928 9956 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10134 8916 10140 8968
rect 10192 8916 10198 8968
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10428 8956 10456 8996
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 12526 9024 12532 9036
rect 11256 8996 12532 9024
rect 10367 8928 10456 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 9968 8888 9996 8916
rect 10226 8888 10232 8900
rect 9968 8860 10232 8888
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 10336 8820 10364 8919
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11256 8965 11284 8996
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 13740 9024 13768 9064
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 14645 9095 14703 9101
rect 14645 9061 14657 9095
rect 14691 9092 14703 9095
rect 14826 9092 14832 9104
rect 14691 9064 14832 9092
rect 14691 9061 14703 9064
rect 14645 9055 14703 9061
rect 14826 9052 14832 9064
rect 14884 9052 14890 9104
rect 13188 8996 13768 9024
rect 14277 9027 14335 9033
rect 11241 8959 11299 8965
rect 10744 8928 10916 8956
rect 10744 8916 10750 8928
rect 10778 8848 10784 8900
rect 10836 8848 10842 8900
rect 10888 8888 10916 8928
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11440 8888 11468 8919
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 11756 8928 12449 8956
rect 11756 8916 11762 8928
rect 12437 8925 12449 8928
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 12618 8916 12624 8968
rect 12676 8916 12682 8968
rect 12894 8916 12900 8968
rect 12952 8916 12958 8968
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8952 13139 8959
rect 13188 8952 13216 8996
rect 14277 8993 14289 9027
rect 14323 9024 14335 9027
rect 14550 9024 14556 9036
rect 14323 8996 14556 9024
rect 14323 8993 14335 8996
rect 14277 8987 14335 8993
rect 13127 8925 13216 8952
rect 13081 8924 13216 8925
rect 13081 8919 13139 8924
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13320 8928 13369 8956
rect 13320 8916 13326 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 13504 8928 13553 8956
rect 13504 8916 13510 8928
rect 13541 8925 13553 8928
rect 13587 8956 13599 8959
rect 14292 8956 14320 8987
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 13587 8928 14320 8956
rect 14461 8959 14519 8965
rect 13587 8925 13599 8928
rect 13541 8919 13599 8925
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 10888 8860 11468 8888
rect 11974 8848 11980 8900
rect 12032 8848 12038 8900
rect 12989 8891 13047 8897
rect 12989 8888 13001 8891
rect 12452 8860 13001 8888
rect 9048 8792 10364 8820
rect 8389 8783 8447 8789
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 10744 8792 10885 8820
rect 10744 8780 10750 8792
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 10873 8783 10931 8789
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 12452 8820 12480 8860
rect 12989 8857 13001 8860
rect 13035 8857 13047 8891
rect 14476 8888 14504 8919
rect 14918 8916 14924 8968
rect 14976 8916 14982 8968
rect 15120 8965 15148 9132
rect 15378 9120 15384 9172
rect 15436 9120 15442 9172
rect 16669 9163 16727 9169
rect 16669 9129 16681 9163
rect 16715 9160 16727 9163
rect 17218 9160 17224 9172
rect 16715 9132 17224 9160
rect 16715 9129 16727 9132
rect 16669 9123 16727 9129
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 15396 9024 15424 9120
rect 15473 9095 15531 9101
rect 15473 9061 15485 9095
rect 15519 9092 15531 9095
rect 15519 9064 15884 9092
rect 15519 9061 15531 9064
rect 15473 9055 15531 9061
rect 15212 8996 15424 9024
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8925 15163 8959
rect 15105 8919 15163 8925
rect 15212 8897 15240 8996
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8956 15347 8959
rect 15378 8956 15384 8968
rect 15335 8928 15384 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 15378 8916 15384 8928
rect 15436 8916 15442 8968
rect 15470 8916 15476 8968
rect 15528 8956 15534 8968
rect 15580 8956 15608 9064
rect 15856 9033 15884 9064
rect 17586 9052 17592 9104
rect 17644 9052 17650 9104
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 8993 15899 9027
rect 17402 9024 17408 9036
rect 15841 8987 15899 8993
rect 16868 8996 17408 9024
rect 15528 8928 15608 8956
rect 16209 8959 16267 8965
rect 15528 8916 15534 8928
rect 16209 8925 16221 8959
rect 16255 8956 16267 8959
rect 16758 8956 16764 8968
rect 16255 8928 16764 8956
rect 16255 8925 16267 8928
rect 16209 8919 16267 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 16868 8965 16896 8996
rect 17402 8984 17408 8996
rect 17460 8984 17466 9036
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 17126 8916 17132 8968
rect 17184 8916 17190 8968
rect 17954 8916 17960 8968
rect 18012 8965 18018 8968
rect 18012 8959 18050 8965
rect 18038 8925 18050 8959
rect 18012 8919 18050 8925
rect 18012 8916 18018 8919
rect 12989 8851 13047 8857
rect 13096 8860 14504 8888
rect 15197 8891 15255 8897
rect 13096 8832 13124 8860
rect 15197 8857 15209 8891
rect 15243 8888 15255 8891
rect 15746 8888 15752 8900
rect 15243 8860 15752 8888
rect 15243 8857 15255 8860
rect 15197 8851 15255 8857
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 17681 8891 17739 8897
rect 17681 8857 17693 8891
rect 17727 8888 17739 8891
rect 18095 8891 18153 8897
rect 18095 8888 18107 8891
rect 17727 8860 18107 8888
rect 17727 8857 17739 8860
rect 17681 8851 17739 8857
rect 18095 8857 18107 8860
rect 18141 8857 18153 8891
rect 18095 8851 18153 8857
rect 11020 8792 12480 8820
rect 11020 8780 11026 8792
rect 13078 8780 13084 8832
rect 13136 8780 13142 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 14274 8820 14280 8832
rect 13412 8792 14280 8820
rect 13412 8780 13418 8792
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 15838 8780 15844 8832
rect 15896 8820 15902 8832
rect 16209 8823 16267 8829
rect 16209 8820 16221 8823
rect 15896 8792 16221 8820
rect 15896 8780 15902 8792
rect 16209 8789 16221 8792
rect 16255 8789 16267 8823
rect 16209 8783 16267 8789
rect 1104 8730 18860 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 16214 8730
rect 16266 8678 16278 8730
rect 16330 8678 16342 8730
rect 16394 8678 16406 8730
rect 16458 8678 16470 8730
rect 16522 8678 18860 8730
rect 1104 8656 18860 8678
rect 6086 8576 6092 8628
rect 6144 8576 6150 8628
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 7558 8616 7564 8628
rect 7340 8588 7564 8616
rect 7340 8576 7346 8588
rect 7558 8576 7564 8588
rect 7616 8616 7622 8628
rect 8757 8619 8815 8625
rect 8757 8616 8769 8619
rect 7616 8588 8769 8616
rect 7616 8576 7622 8588
rect 8757 8585 8769 8588
rect 8803 8585 8815 8619
rect 8757 8579 8815 8585
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 13262 8616 13268 8628
rect 9447 8588 13268 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13817 8619 13875 8625
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 14366 8616 14372 8628
rect 13863 8588 14372 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 15194 8616 15200 8628
rect 14608 8588 15200 8616
rect 14608 8576 14614 8588
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 15838 8576 15844 8628
rect 15896 8576 15902 8628
rect 16942 8616 16948 8628
rect 16040 8588 16948 8616
rect 6454 8548 6460 8560
rect 4172 8520 6460 8548
rect 2038 8440 2044 8492
rect 2096 8440 2102 8492
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 4172 8489 4200 8520
rect 6454 8508 6460 8520
rect 6512 8548 6518 8560
rect 6512 8520 6684 8548
rect 6512 8508 6518 8520
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6178 8480 6184 8492
rect 5767 8452 6184 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6656 8489 6684 8520
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 8018 8548 8024 8560
rect 7064 8520 8024 8548
rect 7064 8508 7070 8520
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 7098 8440 7104 8492
rect 7156 8440 7162 8492
rect 7300 8489 7328 8520
rect 8018 8508 8024 8520
rect 8076 8508 8082 8560
rect 9766 8508 9772 8560
rect 9824 8508 9830 8560
rect 9907 8551 9965 8557
rect 9907 8517 9919 8551
rect 9953 8548 9965 8551
rect 10226 8548 10232 8560
rect 9953 8520 10232 8548
rect 9953 8517 9965 8520
rect 9907 8511 9965 8517
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 12066 8548 12072 8560
rect 10336 8520 12072 8548
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8480 7987 8483
rect 8110 8480 8116 8492
rect 7975 8452 8116 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 3510 8412 3516 8424
rect 2639 8384 3516 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 6420 8384 7420 8412
rect 6420 8372 6426 8384
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 4890 8344 4896 8356
rect 4203 8316 4896 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4890 8304 4896 8316
rect 4948 8304 4954 8356
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 6457 8347 6515 8353
rect 6457 8344 6469 8347
rect 6135 8316 6469 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 6457 8313 6469 8316
rect 6503 8313 6515 8347
rect 6457 8307 6515 8313
rect 7098 8304 7104 8356
rect 7156 8304 7162 8356
rect 7392 8344 7420 8384
rect 7466 8372 7472 8424
rect 7524 8412 7530 8424
rect 7760 8412 7788 8443
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 8570 8440 8576 8492
rect 8628 8480 8634 8492
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8628 8452 8677 8480
rect 8628 8440 8634 8452
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 9306 8480 9312 8492
rect 8895 8452 9312 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9582 8440 9588 8492
rect 9640 8440 9646 8492
rect 9674 8440 9680 8492
rect 9732 8440 9738 8492
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10336 8480 10364 8520
rect 12066 8508 12072 8520
rect 12124 8508 12130 8560
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 13538 8548 13544 8560
rect 12483 8520 13544 8548
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 15856 8548 15884 8576
rect 13648 8520 14688 8548
rect 10100 8452 10364 8480
rect 10100 8440 10106 8452
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11422 8480 11428 8492
rect 11112 8452 11428 8480
rect 11112 8440 11118 8452
rect 11422 8440 11428 8452
rect 11480 8480 11486 8492
rect 11609 8483 11667 8489
rect 11609 8480 11621 8483
rect 11480 8452 11621 8480
rect 11480 8440 11486 8452
rect 11609 8449 11621 8452
rect 11655 8449 11667 8483
rect 11609 8443 11667 8449
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 12710 8480 12716 8492
rect 12575 8452 12716 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 7524 8384 7788 8412
rect 7524 8372 7530 8384
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 9916 8384 11713 8412
rect 9916 8372 9922 8384
rect 11701 8381 11713 8384
rect 11747 8412 11759 8415
rect 11882 8412 11888 8424
rect 11747 8384 11888 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 11882 8372 11888 8384
rect 11940 8412 11946 8424
rect 12360 8412 12388 8443
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 11940 8384 12388 8412
rect 11940 8372 11946 8384
rect 9490 8344 9496 8356
rect 7392 8316 9496 8344
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 10134 8344 10140 8356
rect 10060 8316 10140 8344
rect 2222 8236 2228 8288
rect 2280 8276 2286 8288
rect 8386 8276 8392 8288
rect 2280 8248 8392 8276
rect 2280 8236 2286 8248
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 9766 8276 9772 8306
rect 8628 8254 9772 8276
rect 9824 8254 9830 8306
rect 10060 8294 10088 8316
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 10962 8344 10968 8356
rect 10744 8316 10968 8344
rect 10744 8304 10750 8316
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 12820 8344 12848 8443
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13648 8489 13676 8520
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13412 8452 13645 8480
rect 13412 8440 13418 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 13906 8440 13912 8492
rect 13964 8440 13970 8492
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8480 14427 8483
rect 14458 8480 14464 8492
rect 14415 8452 14464 8480
rect 14415 8449 14427 8452
rect 14369 8443 14427 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14660 8489 14688 8520
rect 15764 8520 15884 8548
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 14844 8412 14872 8443
rect 15470 8440 15476 8492
rect 15528 8440 15534 8492
rect 12943 8384 14136 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 13446 8344 13452 8356
rect 12124 8316 12848 8344
rect 12912 8316 13452 8344
rect 12124 8304 12130 8316
rect 9876 8276 10088 8294
rect 10321 8279 10379 8285
rect 10321 8276 10333 8279
rect 8628 8248 9812 8254
rect 9876 8248 10333 8276
rect 8628 8236 8634 8248
rect 10321 8245 10333 8248
rect 10367 8276 10379 8279
rect 10410 8276 10416 8288
rect 10367 8248 10416 8276
rect 10367 8245 10379 8248
rect 10321 8239 10379 8245
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 12912 8276 12940 8316
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 13633 8347 13691 8353
rect 13633 8313 13645 8347
rect 13679 8344 13691 8347
rect 13814 8344 13820 8356
rect 13679 8316 13820 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 11848 8248 12940 8276
rect 11848 8236 11854 8248
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 13906 8276 13912 8288
rect 13320 8248 13912 8276
rect 13320 8236 13326 8248
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 14108 8276 14136 8384
rect 14660 8384 14872 8412
rect 14274 8304 14280 8356
rect 14332 8304 14338 8356
rect 14660 8344 14688 8384
rect 14384 8316 14688 8344
rect 15764 8344 15792 8520
rect 16040 8480 16068 8588
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17586 8508 17592 8560
rect 17644 8548 17650 8560
rect 17957 8551 18015 8557
rect 17957 8548 17969 8551
rect 17644 8520 17969 8548
rect 17644 8508 17650 8520
rect 17957 8517 17969 8520
rect 18003 8517 18015 8551
rect 17957 8511 18015 8517
rect 15856 8452 16068 8480
rect 16209 8483 16267 8489
rect 15856 8421 15884 8452
rect 16209 8449 16221 8483
rect 16255 8449 16267 8483
rect 16796 8483 16854 8489
rect 16796 8480 16808 8483
rect 16209 8443 16267 8449
rect 16776 8449 16808 8480
rect 16842 8449 16854 8483
rect 16776 8443 16854 8449
rect 15841 8415 15899 8421
rect 15841 8381 15853 8415
rect 15887 8381 15899 8415
rect 16224 8412 16252 8443
rect 16666 8412 16672 8424
rect 16224 8384 16672 8412
rect 15841 8375 15899 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 16776 8344 16804 8443
rect 15764 8316 16804 8344
rect 14384 8276 14412 8316
rect 17770 8304 17776 8356
rect 17828 8344 17834 8356
rect 18141 8347 18199 8353
rect 18141 8344 18153 8347
rect 17828 8316 18153 8344
rect 17828 8304 17834 8316
rect 18141 8313 18153 8316
rect 18187 8313 18199 8347
rect 18141 8307 18199 8313
rect 14108 8248 14412 8276
rect 14642 8236 14648 8288
rect 14700 8236 14706 8288
rect 15930 8236 15936 8288
rect 15988 8276 15994 8288
rect 16301 8279 16359 8285
rect 16301 8276 16313 8279
rect 15988 8248 16313 8276
rect 15988 8236 15994 8248
rect 16301 8245 16313 8248
rect 16347 8245 16359 8279
rect 16301 8239 16359 8245
rect 16574 8236 16580 8288
rect 16632 8276 16638 8288
rect 16899 8279 16957 8285
rect 16899 8276 16911 8279
rect 16632 8248 16911 8276
rect 16632 8236 16638 8248
rect 16899 8245 16911 8248
rect 16945 8245 16957 8279
rect 16899 8239 16957 8245
rect 1104 8186 18860 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 18860 8186
rect 1104 8112 18860 8134
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3602 8072 3608 8084
rect 3467 8044 3608 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 6144 8044 6193 8072
rect 6144 8032 6150 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 11238 8072 11244 8084
rect 9548 8044 11244 8072
rect 9548 8032 9554 8044
rect 11238 8032 11244 8044
rect 11296 8032 11302 8084
rect 12710 8072 12716 8084
rect 11348 8044 12716 8072
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 3016 7908 3525 7936
rect 3016 7896 3022 7908
rect 3513 7905 3525 7908
rect 3559 7905 3571 7939
rect 3620 7936 3648 8032
rect 4709 8007 4767 8013
rect 4709 7973 4721 8007
rect 4755 8004 4767 8007
rect 4890 8004 4896 8016
rect 4755 7976 4896 8004
rect 4755 7973 4767 7976
rect 4709 7967 4767 7973
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 6914 7964 6920 8016
rect 6972 8004 6978 8016
rect 7929 8007 7987 8013
rect 7929 8004 7941 8007
rect 6972 7976 7941 8004
rect 6972 7964 6978 7976
rect 7929 7973 7941 7976
rect 7975 7973 7987 8007
rect 7929 7967 7987 7973
rect 9306 7964 9312 8016
rect 9364 8004 9370 8016
rect 11348 8013 11376 8044
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 11333 8007 11391 8013
rect 11333 8004 11345 8007
rect 9364 7976 11345 8004
rect 9364 7964 9370 7976
rect 11333 7973 11345 7976
rect 11379 7973 11391 8007
rect 11333 7967 11391 7973
rect 12253 8007 12311 8013
rect 12253 7973 12265 8007
rect 12299 8004 12311 8007
rect 12299 7976 12434 8004
rect 12299 7973 12311 7976
rect 12253 7967 12311 7973
rect 4249 7939 4307 7945
rect 4249 7936 4261 7939
rect 3620 7908 4261 7936
rect 3513 7899 3571 7905
rect 4249 7905 4261 7908
rect 4295 7905 4307 7939
rect 4249 7899 4307 7905
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 5534 7936 5540 7948
rect 4847 7908 5540 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7936 6055 7939
rect 6178 7936 6184 7948
rect 6043 7908 6184 7936
rect 6043 7905 6055 7908
rect 5997 7899 6055 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7936 6423 7939
rect 6454 7936 6460 7948
rect 6411 7908 6460 7936
rect 6411 7905 6423 7908
rect 6365 7899 6423 7905
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 7098 7936 7104 7948
rect 6656 7908 7104 7936
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 2314 7828 2320 7880
rect 2372 7828 2378 7880
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2590 7868 2596 7880
rect 2547 7840 2596 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2424 7800 2452 7831
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 3234 7828 3240 7880
rect 3292 7828 3298 7880
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7868 3387 7871
rect 6656 7868 6684 7908
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 8018 7936 8024 7948
rect 7208 7908 8024 7936
rect 3375 7840 6684 7868
rect 6733 7871 6791 7877
rect 3375 7837 3387 7840
rect 3329 7831 3387 7837
rect 6733 7837 6745 7871
rect 6779 7868 6791 7871
rect 7208 7868 7236 7908
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 9950 7936 9956 7948
rect 8352 7908 9956 7936
rect 8352 7896 8358 7908
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10321 7939 10379 7945
rect 10321 7905 10333 7939
rect 10367 7936 10379 7939
rect 10410 7936 10416 7948
rect 10367 7908 10416 7936
rect 10367 7905 10379 7908
rect 10321 7899 10379 7905
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7936 12035 7939
rect 12066 7936 12072 7948
rect 12023 7908 12072 7936
rect 12023 7905 12035 7908
rect 11977 7899 12035 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12406 7936 12434 7976
rect 12894 7964 12900 8016
rect 12952 8004 12958 8016
rect 15289 8007 15347 8013
rect 12952 7976 13584 8004
rect 12952 7964 12958 7976
rect 12406 7908 13492 7936
rect 13464 7880 13492 7908
rect 6779 7840 7236 7868
rect 7285 7871 7343 7877
rect 6779 7837 6791 7840
rect 6733 7831 6791 7837
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 7558 7868 7564 7880
rect 7331 7840 7564 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 3878 7800 3884 7812
rect 2424 7772 3884 7800
rect 3878 7760 3884 7772
rect 3936 7760 3942 7812
rect 6748 7800 6776 7831
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7868 7711 7871
rect 7742 7868 7748 7880
rect 7699 7840 7748 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 6656 7772 6776 7800
rect 7377 7803 7435 7809
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 6656 7732 6684 7772
rect 7377 7769 7389 7803
rect 7423 7800 7435 7803
rect 7944 7800 7972 7831
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 10134 7868 10140 7880
rect 8444 7840 10140 7868
rect 8444 7828 8450 7840
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 10502 7800 10508 7812
rect 7423 7772 10508 7800
rect 7423 7769 7435 7772
rect 7377 7763 7435 7769
rect 10502 7760 10508 7772
rect 10560 7760 10566 7812
rect 11256 7800 11284 7831
rect 11790 7828 11796 7880
rect 11848 7868 11854 7880
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11848 7840 11897 7868
rect 11848 7828 11854 7840
rect 11885 7837 11897 7840
rect 11931 7837 11943 7871
rect 11885 7831 11943 7837
rect 13262 7828 13268 7880
rect 13320 7828 13326 7880
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 13556 7877 13584 7976
rect 15289 7973 15301 8007
rect 15335 8004 15347 8007
rect 15470 8004 15476 8016
rect 15335 7976 15476 8004
rect 15335 7973 15347 7976
rect 15289 7967 15347 7973
rect 15470 7964 15476 7976
rect 15528 8004 15534 8016
rect 15746 8004 15752 8016
rect 15528 7976 15752 8004
rect 15528 7964 15534 7976
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13964 7908 14289 7936
rect 13964 7896 13970 7908
rect 14277 7905 14289 7908
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14734 7896 14740 7948
rect 14792 7896 14798 7948
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 16022 7936 16028 7948
rect 15611 7908 16028 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 13556 7871 13625 7877
rect 13556 7840 13579 7871
rect 13567 7837 13579 7840
rect 13613 7837 13625 7871
rect 13567 7831 13625 7837
rect 13722 7828 13728 7880
rect 13780 7828 13786 7880
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 14642 7868 14648 7880
rect 14424 7840 14648 7868
rect 14424 7828 14430 7840
rect 14642 7828 14648 7840
rect 14700 7828 14706 7880
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 15068 7840 15117 7868
rect 15068 7828 15074 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7868 16543 7871
rect 16574 7868 16580 7880
rect 16531 7840 16580 7868
rect 16531 7837 16543 7840
rect 16485 7831 16543 7837
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 16850 7828 16856 7880
rect 16908 7828 16914 7880
rect 17770 7828 17776 7880
rect 17828 7828 17834 7880
rect 18116 7871 18174 7877
rect 18116 7837 18128 7871
rect 18162 7868 18174 7871
rect 18322 7868 18328 7880
rect 18162 7840 18328 7868
rect 18162 7837 18174 7840
rect 18116 7831 18174 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 12802 7800 12808 7812
rect 11256 7772 12808 7800
rect 12802 7760 12808 7772
rect 12860 7800 12866 7812
rect 13170 7800 13176 7812
rect 12860 7772 13176 7800
rect 12860 7760 12866 7772
rect 13170 7760 13176 7772
rect 13228 7760 13234 7812
rect 13357 7803 13415 7809
rect 13357 7769 13369 7803
rect 13403 7800 13415 7803
rect 14384 7800 14412 7828
rect 13403 7772 14412 7800
rect 13403 7769 13415 7772
rect 13357 7763 13415 7769
rect 16206 7760 16212 7812
rect 16264 7760 16270 7812
rect 16942 7760 16948 7812
rect 17000 7800 17006 7812
rect 17497 7803 17555 7809
rect 17497 7800 17509 7803
rect 17000 7772 17509 7800
rect 17000 7760 17006 7772
rect 17497 7769 17509 7772
rect 17543 7769 17555 7803
rect 17497 7763 17555 7769
rect 2087 7704 6684 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6788 7704 6929 7732
rect 6788 7692 6794 7704
rect 6917 7701 6929 7704
rect 6963 7701 6975 7735
rect 6917 7695 6975 7701
rect 7466 7692 7472 7744
rect 7524 7692 7530 7744
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 7834 7732 7840 7744
rect 7699 7704 7840 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 9732 7704 10609 7732
rect 9732 7692 9738 7704
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10597 7695 10655 7701
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 13081 7735 13139 7741
rect 13081 7732 13093 7735
rect 12768 7704 13093 7732
rect 12768 7692 12774 7704
rect 13081 7701 13093 7704
rect 13127 7701 13139 7735
rect 13081 7695 13139 7701
rect 18138 7692 18144 7744
rect 18196 7741 18202 7744
rect 18196 7735 18245 7741
rect 18196 7701 18199 7735
rect 18233 7701 18245 7735
rect 18196 7695 18245 7701
rect 18196 7692 18202 7695
rect 1104 7642 18860 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 16214 7642
rect 16266 7590 16278 7642
rect 16330 7590 16342 7642
rect 16394 7590 16406 7642
rect 16458 7590 16470 7642
rect 16522 7590 18860 7642
rect 1104 7568 18860 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 2740 7500 5733 7528
rect 2740 7488 2746 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 6851 7531 6909 7537
rect 6851 7497 6863 7531
rect 6897 7528 6909 7531
rect 8110 7528 8116 7540
rect 6897 7500 8116 7528
rect 6897 7497 6909 7500
rect 6851 7491 6909 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7528 8999 7531
rect 10226 7528 10232 7540
rect 8987 7500 10232 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11020 7500 13216 7528
rect 11020 7488 11026 7500
rect 5000 7432 5856 7460
rect 5000 7404 5028 7432
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2130 7392 2136 7404
rect 1903 7364 2136 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2406 7352 2412 7404
rect 2464 7352 2470 7404
rect 2498 7352 2504 7404
rect 2556 7352 2562 7404
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2682 7392 2688 7404
rect 2639 7364 2688 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 2792 7324 2820 7355
rect 3234 7352 3240 7404
rect 3292 7352 3298 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5828 7401 5856 7432
rect 6362 7420 6368 7472
rect 6420 7460 6426 7472
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 6420 7432 6653 7460
rect 6420 7420 6426 7432
rect 6641 7429 6653 7432
rect 6687 7460 6699 7463
rect 6730 7460 6736 7472
rect 6687 7432 6736 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 6730 7420 6736 7432
rect 6788 7460 6794 7472
rect 8128 7460 8156 7488
rect 9582 7460 9588 7472
rect 6788 7432 7788 7460
rect 8128 7432 9588 7460
rect 6788 7420 6794 7432
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 1811 7296 2820 7324
rect 3053 7327 3111 7333
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 3053 7293 3065 7327
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 2372 7228 2728 7256
rect 2372 7216 2378 7228
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 2590 7188 2596 7200
rect 2179 7160 2596 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 2700 7188 2728 7228
rect 2774 7216 2780 7268
rect 2832 7256 2838 7268
rect 3068 7256 3096 7287
rect 2832 7228 3096 7256
rect 3252 7256 3280 7352
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4856 7296 4905 7324
rect 4856 7284 4862 7296
rect 4893 7293 4905 7296
rect 4939 7324 4951 7327
rect 5644 7324 5672 7355
rect 4939 7296 5672 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 5353 7259 5411 7265
rect 5353 7256 5365 7259
rect 3252 7228 5365 7256
rect 2832 7216 2838 7228
rect 5353 7225 5365 7228
rect 5399 7225 5411 7259
rect 7098 7256 7104 7268
rect 5353 7219 5411 7225
rect 6840 7228 7104 7256
rect 6840 7197 6868 7228
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 7668 7256 7696 7355
rect 7760 7333 7788 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 10410 7420 10416 7472
rect 10468 7460 10474 7472
rect 13188 7460 13216 7500
rect 13354 7488 13360 7540
rect 13412 7488 13418 7540
rect 16758 7488 16764 7540
rect 16816 7488 16822 7540
rect 13722 7460 13728 7472
rect 10468 7432 12020 7460
rect 10468 7420 10474 7432
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8110 7392 8116 7404
rect 7975 7364 8116 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 8570 7352 8576 7404
rect 8628 7352 8634 7404
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9364 7364 10333 7392
rect 9364 7352 9370 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 11882 7352 11888 7404
rect 11940 7352 11946 7404
rect 11992 7401 12020 7432
rect 13188 7432 13728 7460
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 12066 7352 12072 7404
rect 12124 7352 12130 7404
rect 13188 7401 13216 7432
rect 13722 7420 13728 7432
rect 13780 7420 13786 7472
rect 15470 7460 15476 7472
rect 15120 7432 15476 7460
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7324 7803 7327
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 7791 7296 8677 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 8665 7293 8677 7296
rect 8711 7324 8723 7327
rect 10042 7324 10048 7336
rect 8711 7296 10048 7324
rect 8711 7293 8723 7296
rect 8665 7287 8723 7293
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 10413 7327 10471 7333
rect 10413 7293 10425 7327
rect 10459 7324 10471 7327
rect 11609 7327 11667 7333
rect 11609 7324 11621 7327
rect 10459 7296 11621 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 11609 7293 11621 7296
rect 11655 7293 11667 7327
rect 11609 7287 11667 7293
rect 8754 7256 8760 7268
rect 7668 7228 8760 7256
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 10689 7259 10747 7265
rect 10689 7225 10701 7259
rect 10735 7256 10747 7259
rect 11882 7256 11888 7268
rect 10735 7228 11888 7256
rect 10735 7225 10747 7228
rect 10689 7219 10747 7225
rect 11882 7216 11888 7228
rect 11940 7216 11946 7268
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 2700 7160 3433 7188
rect 3421 7157 3433 7160
rect 3467 7157 3479 7191
rect 3421 7151 3479 7157
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 7006 7148 7012 7200
rect 7064 7148 7070 7200
rect 7469 7191 7527 7197
rect 7469 7157 7481 7191
rect 7515 7188 7527 7191
rect 8478 7188 8484 7200
rect 7515 7160 8484 7188
rect 7515 7157 7527 7160
rect 7469 7151 7527 7157
rect 8478 7148 8484 7160
rect 8536 7188 8542 7200
rect 12268 7188 12296 7355
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 15120 7401 15148 7432
rect 15470 7420 15476 7432
rect 15528 7420 15534 7472
rect 15930 7420 15936 7472
rect 15988 7420 15994 7472
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13504 7364 13921 7392
rect 13504 7352 13510 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7361 15163 7395
rect 15105 7355 15163 7361
rect 15286 7352 15292 7404
rect 15344 7352 15350 7404
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16022 7392 16028 7404
rect 15795 7364 16028 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 17000 7364 17877 7392
rect 17000 7352 17006 7364
rect 17865 7361 17877 7364
rect 17911 7361 17923 7395
rect 17865 7355 17923 7361
rect 18138 7352 18144 7404
rect 18196 7352 18202 7404
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 13262 7324 13268 7336
rect 13044 7296 13268 7324
rect 13044 7284 13050 7296
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 13814 7284 13820 7336
rect 13872 7284 13878 7336
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17221 7327 17279 7333
rect 17221 7324 17233 7327
rect 16908 7296 17233 7324
rect 16908 7284 16914 7296
rect 17221 7293 17233 7296
rect 17267 7293 17279 7327
rect 17221 7287 17279 7293
rect 14274 7216 14280 7268
rect 14332 7216 14338 7268
rect 15102 7216 15108 7268
rect 15160 7216 15166 7268
rect 8536 7160 12296 7188
rect 8536 7148 8542 7160
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16117 7191 16175 7197
rect 16117 7188 16129 7191
rect 15804 7160 16129 7188
rect 15804 7148 15810 7160
rect 16117 7157 16129 7160
rect 16163 7157 16175 7191
rect 16117 7151 16175 7157
rect 1104 7098 18860 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 18860 7098
rect 1104 7024 18860 7046
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 2774 6984 2780 6996
rect 2464 6956 2780 6984
rect 2464 6944 2470 6956
rect 2774 6944 2780 6956
rect 2832 6944 2838 6996
rect 3418 6984 3424 6996
rect 2884 6956 3424 6984
rect 1670 6876 1676 6928
rect 1728 6916 1734 6928
rect 2884 6916 2912 6956
rect 3418 6944 3424 6956
rect 3476 6984 3482 6996
rect 4062 6984 4068 6996
rect 3476 6956 4068 6984
rect 3476 6944 3482 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 4982 6984 4988 6996
rect 4571 6956 4988 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 7929 6987 7987 6993
rect 7929 6953 7941 6987
rect 7975 6984 7987 6987
rect 17034 6984 17040 6996
rect 7975 6956 17040 6984
rect 7975 6953 7987 6956
rect 7929 6947 7987 6953
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 1728 6888 2912 6916
rect 2976 6888 6960 6916
rect 1728 6876 1734 6888
rect 2869 6851 2927 6857
rect 2869 6817 2881 6851
rect 2915 6848 2927 6851
rect 2976 6848 3004 6888
rect 2915 6820 3004 6848
rect 2915 6817 2927 6820
rect 2869 6811 2927 6817
rect 4246 6808 4252 6860
rect 4304 6808 4310 6860
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 2314 6740 2320 6792
rect 2372 6780 2378 6792
rect 2409 6783 2467 6789
rect 2409 6780 2421 6783
rect 2372 6752 2421 6780
rect 2372 6740 2378 6752
rect 2409 6749 2421 6752
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 2498 6740 2504 6792
rect 2556 6740 2562 6792
rect 2590 6740 2596 6792
rect 2648 6740 2654 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 2685 6715 2743 6721
rect 2685 6681 2697 6715
rect 2731 6712 2743 6715
rect 2866 6712 2872 6724
rect 2731 6684 2872 6712
rect 2731 6681 2743 6684
rect 2685 6675 2743 6681
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 3602 6644 3608 6656
rect 2188 6616 3608 6644
rect 2188 6604 2194 6616
rect 3602 6604 3608 6616
rect 3660 6644 3666 6656
rect 4172 6644 4200 6743
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 6472 6780 6500 6811
rect 6730 6808 6736 6860
rect 6788 6808 6794 6860
rect 6822 6780 6828 6792
rect 6472 6752 6828 6780
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 6932 6712 6960 6888
rect 7006 6876 7012 6928
rect 7064 6916 7070 6928
rect 7561 6919 7619 6925
rect 7561 6916 7573 6919
rect 7064 6888 7573 6916
rect 7064 6876 7070 6888
rect 7561 6885 7573 6888
rect 7607 6885 7619 6919
rect 7561 6879 7619 6885
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 9861 6919 9919 6925
rect 9861 6916 9873 6919
rect 8168 6888 9873 6916
rect 8168 6876 8174 6888
rect 9861 6885 9873 6888
rect 9907 6885 9919 6919
rect 9861 6879 9919 6885
rect 10612 6888 10824 6916
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 10612 6848 10640 6888
rect 10796 6857 10824 6888
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 13078 6916 13084 6928
rect 10928 6888 13084 6916
rect 10928 6876 10934 6888
rect 9640 6820 10640 6848
rect 10781 6851 10839 6857
rect 9640 6808 9646 6820
rect 10781 6817 10793 6851
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11072 6848 11284 6856
rect 11425 6851 11483 6857
rect 11425 6848 11437 6851
rect 11020 6828 11437 6848
rect 11020 6820 11100 6828
rect 11256 6820 11437 6828
rect 11020 6808 11026 6820
rect 11425 6817 11437 6820
rect 11471 6817 11483 6851
rect 11425 6811 11483 6817
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 9490 6783 9548 6789
rect 9490 6749 9502 6783
rect 9536 6749 9548 6783
rect 9490 6743 9548 6749
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6780 10011 6783
rect 11054 6780 11060 6792
rect 9999 6752 11060 6780
rect 9999 6749 10011 6752
rect 9953 6743 10011 6749
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 6932 6684 7941 6712
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 7929 6675 7987 6681
rect 8665 6715 8723 6721
rect 8665 6681 8677 6715
rect 8711 6712 8723 6715
rect 8754 6712 8760 6724
rect 8711 6684 8760 6712
rect 8711 6681 8723 6684
rect 8665 6675 8723 6681
rect 8754 6672 8760 6684
rect 8812 6712 8818 6724
rect 9505 6712 9533 6743
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11532 6789 11560 6888
rect 13078 6876 13084 6888
rect 13136 6916 13142 6928
rect 13449 6919 13507 6925
rect 13449 6916 13461 6919
rect 13136 6888 13461 6916
rect 13136 6876 13142 6888
rect 13449 6885 13461 6888
rect 13495 6885 13507 6919
rect 13449 6879 13507 6885
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6848 13047 6851
rect 13035 6820 13400 6848
rect 13035 6817 13047 6820
rect 12989 6811 13047 6817
rect 13372 6792 13400 6820
rect 14274 6808 14280 6860
rect 14332 6848 14338 6860
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 14332 6820 14657 6848
rect 14332 6808 14338 6820
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 14645 6811 14703 6817
rect 14826 6808 14832 6860
rect 14884 6808 14890 6860
rect 16945 6851 17003 6857
rect 16945 6848 16957 6851
rect 15488 6820 16957 6848
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 12710 6740 12716 6792
rect 12768 6740 12774 6792
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6780 12863 6783
rect 12894 6780 12900 6792
rect 12851 6752 12900 6780
rect 12851 6749 12863 6752
rect 12805 6743 12863 6749
rect 10042 6712 10048 6724
rect 8812 6684 10048 6712
rect 8812 6672 8818 6684
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 12066 6712 12072 6724
rect 10336 6684 12072 6712
rect 8018 6644 8024 6656
rect 3660 6616 8024 6644
rect 3660 6604 3666 6616
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 9306 6604 9312 6656
rect 9364 6604 9370 6656
rect 9493 6647 9551 6653
rect 9493 6613 9505 6647
rect 9539 6644 9551 6647
rect 9674 6644 9680 6656
rect 9539 6616 9680 6644
rect 9539 6613 9551 6616
rect 9493 6607 9551 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10336 6653 10364 6684
rect 12066 6672 12072 6684
rect 12124 6672 12130 6724
rect 12820 6712 12848 6743
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 12406 6684 12848 6712
rect 13280 6712 13308 6743
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 14844 6780 14872 6808
rect 13412 6752 14872 6780
rect 13412 6740 13418 6752
rect 15194 6740 15200 6792
rect 15252 6740 15258 6792
rect 15488 6724 15516 6820
rect 16945 6817 16957 6820
rect 16991 6817 17003 6851
rect 16945 6811 17003 6817
rect 15746 6740 15752 6792
rect 15804 6740 15810 6792
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 16172 6752 16405 6780
rect 16172 6740 16178 6752
rect 16393 6749 16405 6752
rect 16439 6780 16451 6783
rect 16574 6780 16580 6792
rect 16439 6752 16580 6780
rect 16439 6749 16451 6752
rect 16393 6743 16451 6749
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6780 16727 6783
rect 16850 6780 16856 6792
rect 16715 6752 16856 6780
rect 16715 6749 16727 6752
rect 16669 6743 16727 6749
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 15470 6712 15476 6724
rect 13280 6684 15476 6712
rect 10321 6647 10379 6653
rect 10321 6613 10333 6647
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 10689 6647 10747 6653
rect 10689 6613 10701 6647
rect 10735 6644 10747 6647
rect 11054 6644 11060 6656
rect 10735 6616 11060 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11885 6647 11943 6653
rect 11885 6613 11897 6647
rect 11931 6644 11943 6647
rect 12406 6644 12434 6684
rect 15470 6672 15476 6684
rect 15528 6672 15534 6724
rect 11931 6616 12434 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 12989 6647 13047 6653
rect 12989 6644 13001 6647
rect 12860 6616 13001 6644
rect 12860 6604 12866 6616
rect 12989 6613 13001 6616
rect 13035 6613 13047 6647
rect 12989 6607 13047 6613
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 14458 6644 14464 6656
rect 14231 6616 14464 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 14550 6604 14556 6656
rect 14608 6604 14614 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 15381 6647 15439 6653
rect 15381 6644 15393 6647
rect 14700 6616 15393 6644
rect 14700 6604 14706 6616
rect 15381 6613 15393 6616
rect 15427 6613 15439 6647
rect 15381 6607 15439 6613
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15746 6644 15752 6656
rect 15620 6616 15752 6644
rect 15620 6604 15626 6616
rect 15746 6604 15752 6616
rect 15804 6644 15810 6656
rect 17236 6644 17264 6743
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17368 6752 18061 6780
rect 17368 6740 17374 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18414 6740 18420 6792
rect 18472 6740 18478 6792
rect 15804 6616 17264 6644
rect 15804 6604 15810 6616
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 18417 6647 18475 6653
rect 18417 6644 18429 6647
rect 18380 6616 18429 6644
rect 18380 6604 18386 6616
rect 18417 6613 18429 6616
rect 18463 6613 18475 6647
rect 18417 6607 18475 6613
rect 1104 6554 18860 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 16214 6554
rect 16266 6502 16278 6554
rect 16330 6502 16342 6554
rect 16394 6502 16406 6554
rect 16458 6502 16470 6554
rect 16522 6502 18860 6554
rect 1104 6480 18860 6502
rect 1857 6443 1915 6449
rect 1857 6409 1869 6443
rect 1903 6440 1915 6443
rect 2222 6440 2228 6452
rect 1903 6412 2228 6440
rect 1903 6409 1915 6412
rect 1857 6403 1915 6409
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2961 6443 3019 6449
rect 2961 6440 2973 6443
rect 2556 6412 2973 6440
rect 2556 6400 2562 6412
rect 2961 6409 2973 6412
rect 3007 6409 3019 6443
rect 2961 6403 3019 6409
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 3292 6412 4568 6440
rect 3292 6400 3298 6412
rect 2317 6375 2375 6381
rect 2317 6341 2329 6375
rect 2363 6372 2375 6375
rect 2406 6372 2412 6384
rect 2363 6344 2412 6372
rect 2363 6341 2375 6344
rect 2317 6335 2375 6341
rect 2406 6332 2412 6344
rect 2464 6372 2470 6384
rect 2464 6344 4108 6372
rect 2464 6332 2470 6344
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1820 6276 2145 6304
rect 1820 6264 1826 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2222 6264 2228 6316
rect 2280 6264 2286 6316
rect 3234 6304 3240 6316
rect 2746 6276 3240 6304
rect 1854 6196 1860 6248
rect 1912 6236 1918 6248
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 1912 6208 2605 6236
rect 1912 6196 1918 6208
rect 2593 6205 2605 6208
rect 2639 6236 2651 6239
rect 2746 6236 2774 6276
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3326 6264 3332 6316
rect 3384 6264 3390 6316
rect 3436 6313 3464 6344
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 2639 6208 2774 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 3620 6168 3648 6267
rect 3878 6264 3884 6316
rect 3936 6264 3942 6316
rect 4080 6313 4108 6344
rect 4540 6313 4568 6412
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 6788 6412 7849 6440
rect 6788 6400 6794 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 9953 6443 10011 6449
rect 9953 6409 9965 6443
rect 9999 6440 10011 6443
rect 10502 6440 10508 6452
rect 9999 6412 10508 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10836 6412 10977 6440
rect 10836 6400 10842 6412
rect 10965 6409 10977 6412
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 14734 6440 14740 6452
rect 14599 6412 14740 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 16301 6443 16359 6449
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 17310 6440 17316 6452
rect 16347 6412 17316 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 5920 6344 6684 6372
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 4356 6168 4384 6267
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 5920 6313 5948 6344
rect 6656 6316 6684 6344
rect 8588 6344 9628 6372
rect 8588 6316 8616 6344
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 4948 6276 4997 6304
rect 4948 6264 4954 6276
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6304 6147 6307
rect 6135 6276 6592 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 5184 6168 5212 6267
rect 6564 6245 6592 6276
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6696 6276 6745 6304
rect 6696 6264 6702 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6304 7803 6307
rect 8570 6304 8576 6316
rect 7791 6276 8576 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 9600 6313 9628 6344
rect 10042 6332 10048 6384
rect 10100 6372 10106 6384
rect 10100 6344 11008 6372
rect 10100 6332 10106 6344
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 9858 6304 9864 6316
rect 9815 6276 9864 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 6549 6239 6607 6245
rect 6549 6205 6561 6239
rect 6595 6236 6607 6239
rect 8021 6239 8079 6245
rect 6595 6208 6776 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 6748 6180 6776 6208
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 2280 6140 3648 6168
rect 3712 6140 4384 6168
rect 4448 6140 5212 6168
rect 2280 6128 2286 6140
rect 2501 6103 2559 6109
rect 2501 6069 2513 6103
rect 2547 6100 2559 6103
rect 3326 6100 3332 6112
rect 2547 6072 3332 6100
rect 2547 6069 2559 6072
rect 2501 6063 2559 6069
rect 3326 6060 3332 6072
rect 3384 6100 3390 6112
rect 3712 6100 3740 6140
rect 3384 6072 3740 6100
rect 3384 6060 3390 6072
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4448 6100 4476 6140
rect 6730 6128 6736 6180
rect 6788 6128 6794 6180
rect 8036 6168 8064 6199
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8168 6208 9045 6236
rect 8168 6196 8174 6208
rect 9033 6205 9045 6208
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9784 6236 9812 6267
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 10192 6276 10425 6304
rect 10192 6264 10198 6276
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 10888 6236 10916 6267
rect 9171 6208 9812 6236
rect 10244 6208 10916 6236
rect 10980 6236 11008 6344
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 14461 6375 14519 6381
rect 14461 6372 14473 6375
rect 13320 6344 14473 6372
rect 13320 6332 13326 6344
rect 14461 6341 14473 6344
rect 14507 6372 14519 6375
rect 14642 6372 14648 6384
rect 14507 6344 14648 6372
rect 14507 6341 14519 6344
rect 14461 6335 14519 6341
rect 14642 6332 14648 6344
rect 14700 6332 14706 6384
rect 15102 6332 15108 6384
rect 15160 6372 15166 6384
rect 15933 6375 15991 6381
rect 15933 6372 15945 6375
rect 15160 6344 15945 6372
rect 15160 6332 15166 6344
rect 15933 6341 15945 6344
rect 15979 6341 15991 6375
rect 15933 6335 15991 6341
rect 17681 6375 17739 6381
rect 17681 6341 17693 6375
rect 17727 6372 17739 6375
rect 17770 6372 17776 6384
rect 17727 6344 17776 6372
rect 17727 6341 17739 6344
rect 17681 6335 17739 6341
rect 17770 6332 17776 6344
rect 17828 6332 17834 6384
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11609 6307 11667 6313
rect 11609 6304 11621 6307
rect 11296 6276 11621 6304
rect 11296 6264 11302 6276
rect 11609 6273 11621 6276
rect 11655 6273 11667 6307
rect 11609 6267 11667 6273
rect 12710 6264 12716 6316
rect 12768 6264 12774 6316
rect 12802 6264 12808 6316
rect 12860 6264 12866 6316
rect 13078 6264 13084 6316
rect 13136 6264 13142 6316
rect 15746 6264 15752 6316
rect 15804 6264 15810 6316
rect 16022 6264 16028 6316
rect 16080 6264 16086 6316
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 10980 6208 13001 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 8754 6168 8760 6180
rect 8036 6140 8760 6168
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 9582 6128 9588 6180
rect 9640 6168 9646 6180
rect 10244 6168 10272 6208
rect 12989 6205 13001 6208
rect 13035 6236 13047 6239
rect 13354 6236 13360 6248
rect 13035 6208 13360 6236
rect 13035 6205 13047 6208
rect 12989 6199 13047 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6236 14795 6239
rect 14826 6236 14832 6248
rect 14783 6208 14832 6236
rect 14783 6205 14795 6208
rect 14737 6199 14795 6205
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 16132 6236 16160 6267
rect 17310 6264 17316 6316
rect 17368 6264 17374 6316
rect 15948 6208 16160 6236
rect 15948 6180 15976 6208
rect 9640 6140 10272 6168
rect 9640 6128 9646 6140
rect 10318 6128 10324 6180
rect 10376 6168 10382 6180
rect 10597 6171 10655 6177
rect 10597 6168 10609 6171
rect 10376 6140 10609 6168
rect 10376 6128 10382 6140
rect 10597 6137 10609 6140
rect 10643 6168 10655 6171
rect 12529 6171 12587 6177
rect 10643 6140 12434 6168
rect 10643 6137 10655 6140
rect 10597 6131 10655 6137
rect 4028 6072 4476 6100
rect 4028 6060 4034 6072
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 5077 6103 5135 6109
rect 5077 6100 5089 6103
rect 4672 6072 5089 6100
rect 4672 6060 4678 6072
rect 5077 6069 5089 6072
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 5500 6072 5917 6100
rect 5500 6060 5506 6072
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6144 6072 6929 6100
rect 6144 6060 6150 6072
rect 6917 6069 6929 6072
rect 6963 6069 6975 6103
rect 6917 6063 6975 6069
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 7377 6103 7435 6109
rect 7377 6100 7389 6103
rect 7156 6072 7389 6100
rect 7156 6060 7162 6072
rect 7377 6069 7389 6072
rect 7423 6069 7435 6103
rect 7377 6063 7435 6069
rect 8662 6060 8668 6112
rect 8720 6060 8726 6112
rect 11790 6060 11796 6112
rect 11848 6060 11854 6112
rect 12406 6100 12434 6140
rect 12529 6137 12541 6171
rect 12575 6168 12587 6171
rect 13998 6168 14004 6180
rect 12575 6140 14004 6168
rect 12575 6137 12587 6140
rect 12529 6131 12587 6137
rect 13998 6128 14004 6140
rect 14056 6128 14062 6180
rect 15930 6128 15936 6180
rect 15988 6128 15994 6180
rect 17681 6171 17739 6177
rect 17681 6137 17693 6171
rect 17727 6168 17739 6171
rect 18322 6168 18328 6180
rect 17727 6140 18328 6168
rect 17727 6137 17739 6140
rect 17681 6131 17739 6137
rect 18322 6128 18328 6140
rect 18380 6128 18386 6180
rect 12986 6100 12992 6112
rect 12406 6072 12992 6100
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13906 6060 13912 6112
rect 13964 6060 13970 6112
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14366 6100 14372 6112
rect 14139 6072 14372 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 1104 6010 18860 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 18860 6010
rect 1104 5936 18860 5958
rect 2406 5856 2412 5908
rect 2464 5856 2470 5908
rect 4157 5899 4215 5905
rect 4157 5865 4169 5899
rect 4203 5896 4215 5899
rect 4430 5896 4436 5908
rect 4203 5868 4436 5896
rect 4203 5865 4215 5868
rect 4157 5859 4215 5865
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4617 5899 4675 5905
rect 4617 5865 4629 5899
rect 4663 5896 4675 5899
rect 4798 5896 4804 5908
rect 4663 5868 4804 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 9769 5899 9827 5905
rect 9769 5896 9781 5899
rect 9640 5868 9781 5896
rect 9640 5856 9646 5868
rect 9769 5865 9781 5868
rect 9815 5865 9827 5899
rect 9769 5859 9827 5865
rect 12710 5856 12716 5908
rect 12768 5896 12774 5908
rect 12897 5899 12955 5905
rect 12897 5896 12909 5899
rect 12768 5868 12909 5896
rect 12768 5856 12774 5868
rect 12897 5865 12909 5868
rect 12943 5865 12955 5899
rect 12897 5859 12955 5865
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 13817 5899 13875 5905
rect 13817 5896 13829 5899
rect 13412 5868 13829 5896
rect 13412 5856 13418 5868
rect 13817 5865 13829 5868
rect 13863 5896 13875 5899
rect 16022 5896 16028 5908
rect 13863 5868 16028 5896
rect 13863 5865 13875 5868
rect 13817 5859 13875 5865
rect 16022 5856 16028 5868
rect 16080 5856 16086 5908
rect 17957 5899 18015 5905
rect 17957 5865 17969 5899
rect 18003 5896 18015 5899
rect 18414 5896 18420 5908
rect 18003 5868 18420 5896
rect 18003 5865 18015 5868
rect 17957 5859 18015 5865
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 3326 5788 3332 5840
rect 3384 5828 3390 5840
rect 4341 5831 4399 5837
rect 4341 5828 4353 5831
rect 3384 5800 4353 5828
rect 3384 5788 3390 5800
rect 4341 5797 4353 5800
rect 4387 5797 4399 5831
rect 5350 5828 5356 5840
rect 4341 5791 4399 5797
rect 4908 5800 5356 5828
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5760 2835 5763
rect 3142 5760 3148 5772
rect 2823 5732 3148 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 4908 5769 4936 5800
rect 5350 5788 5356 5800
rect 5408 5788 5414 5840
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 3988 5732 4905 5760
rect 1854 5652 1860 5704
rect 1912 5652 1918 5704
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 1995 5664 2605 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 2958 5692 2964 5704
rect 2915 5664 2964 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 2700 5624 2728 5655
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3050 5652 3056 5704
rect 3108 5652 3114 5704
rect 3326 5624 3332 5636
rect 2700 5596 3332 5624
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 3988 5633 4016 5732
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 6086 5760 6092 5772
rect 5123 5732 6092 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 7098 5720 7104 5772
rect 7156 5720 7162 5772
rect 8588 5760 8616 5856
rect 11974 5760 11980 5772
rect 8588 5732 9996 5760
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4488 5664 4813 5692
rect 4488 5652 4494 5664
rect 4801 5661 4813 5664
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 3973 5627 4031 5633
rect 3973 5593 3985 5627
rect 4019 5593 4031 5627
rect 3973 5587 4031 5593
rect 4189 5627 4247 5633
rect 4189 5593 4201 5627
rect 4235 5624 4247 5627
rect 4816 5624 4844 5655
rect 4982 5652 4988 5704
rect 5040 5652 5046 5704
rect 5442 5652 5448 5704
rect 5500 5652 5506 5704
rect 5599 5695 5657 5701
rect 5599 5661 5611 5695
rect 5645 5692 5657 5695
rect 5994 5692 6000 5704
rect 5645 5664 6000 5692
rect 5645 5661 5657 5664
rect 5599 5655 5657 5661
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6822 5652 6828 5704
rect 6880 5652 6886 5704
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 9180 5664 9321 5692
rect 9180 5652 9186 5664
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5692 9827 5695
rect 9858 5692 9864 5704
rect 9815 5664 9864 5692
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 5074 5624 5080 5636
rect 4235 5596 4752 5624
rect 4816 5596 5080 5624
rect 4235 5593 4247 5596
rect 4189 5587 4247 5593
rect 4724 5568 4752 5596
rect 5074 5584 5080 5596
rect 5132 5584 5138 5636
rect 8110 5584 8116 5636
rect 8168 5584 8174 5636
rect 9508 5624 9536 5655
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 9968 5701 9996 5732
rect 10520 5732 11980 5760
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10318 5652 10324 5704
rect 10376 5652 10382 5704
rect 10520 5633 10548 5732
rect 11974 5720 11980 5732
rect 12032 5760 12038 5772
rect 12032 5732 13676 5760
rect 12032 5720 12038 5732
rect 11790 5652 11796 5704
rect 11848 5652 11854 5704
rect 12618 5652 12624 5704
rect 12676 5652 12682 5704
rect 12713 5695 12771 5701
rect 12713 5661 12725 5695
rect 12759 5692 12771 5695
rect 12894 5692 12900 5704
rect 12759 5664 12900 5692
rect 12759 5661 12771 5664
rect 12713 5655 12771 5661
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 13078 5652 13084 5704
rect 13136 5692 13142 5704
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 13136 5664 13185 5692
rect 13136 5652 13142 5664
rect 13173 5661 13185 5664
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13354 5652 13360 5704
rect 13412 5652 13418 5704
rect 13648 5701 13676 5732
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 14185 5763 14243 5769
rect 14185 5760 14197 5763
rect 13964 5732 14197 5760
rect 13964 5720 13970 5732
rect 14185 5729 14197 5732
rect 14231 5729 14243 5763
rect 14185 5723 14243 5729
rect 14458 5720 14464 5772
rect 14516 5720 14522 5772
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 15933 5763 15991 5769
rect 15933 5760 15945 5763
rect 14608 5732 15945 5760
rect 14608 5720 14614 5732
rect 15933 5729 15945 5732
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 16114 5720 16120 5772
rect 16172 5760 16178 5772
rect 16393 5763 16451 5769
rect 16393 5760 16405 5763
rect 16172 5732 16405 5760
rect 16172 5720 16178 5732
rect 16393 5729 16405 5732
rect 16439 5729 16451 5763
rect 16393 5723 16451 5729
rect 16574 5720 16580 5772
rect 16632 5760 16638 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 16632 5732 17049 5760
rect 16632 5720 16638 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 17218 5652 17224 5704
rect 17276 5652 17282 5704
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 18141 5695 18199 5701
rect 18141 5692 18153 5695
rect 17828 5664 18153 5692
rect 17828 5652 17834 5664
rect 18141 5661 18153 5664
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 10505 5627 10563 5633
rect 10505 5624 10517 5627
rect 9508 5596 10517 5624
rect 10505 5593 10517 5596
rect 10551 5593 10563 5627
rect 10505 5587 10563 5593
rect 11606 5584 11612 5636
rect 11664 5624 11670 5636
rect 11885 5627 11943 5633
rect 11885 5624 11897 5627
rect 11664 5596 11897 5624
rect 11664 5584 11670 5596
rect 11885 5593 11897 5596
rect 11931 5593 11943 5627
rect 11885 5587 11943 5593
rect 13265 5627 13323 5633
rect 13265 5593 13277 5627
rect 13311 5624 13323 5627
rect 14090 5624 14096 5636
rect 13311 5596 14096 5624
rect 13311 5593 13323 5596
rect 13265 5587 13323 5593
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 16850 5624 16856 5636
rect 15686 5596 16856 5624
rect 16850 5584 16856 5596
rect 16908 5584 16914 5636
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 5813 5559 5871 5565
rect 5813 5556 5825 5559
rect 4764 5528 5825 5556
rect 4764 5516 4770 5528
rect 5813 5525 5825 5528
rect 5859 5525 5871 5559
rect 5813 5519 5871 5525
rect 8938 5516 8944 5568
rect 8996 5516 9002 5568
rect 9401 5559 9459 5565
rect 9401 5525 9413 5559
rect 9447 5556 9459 5559
rect 9674 5556 9680 5568
rect 9447 5528 9680 5556
rect 9447 5525 9459 5528
rect 9401 5519 9459 5525
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 1104 5466 18860 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 16214 5466
rect 16266 5414 16278 5466
rect 16330 5414 16342 5466
rect 16394 5414 16406 5466
rect 16458 5414 16470 5466
rect 16522 5414 18860 5466
rect 1104 5392 18860 5414
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 2317 5355 2375 5361
rect 2317 5352 2329 5355
rect 2280 5324 2329 5352
rect 2280 5312 2286 5324
rect 2317 5321 2329 5324
rect 2363 5321 2375 5355
rect 2317 5315 2375 5321
rect 3234 5312 3240 5364
rect 3292 5312 3298 5364
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4479 5324 4936 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 1719 5256 2452 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 2424 5225 2452 5256
rect 4706 5244 4712 5296
rect 4764 5244 4770 5296
rect 4798 5244 4804 5296
rect 4856 5284 4862 5296
rect 4908 5284 4936 5324
rect 4982 5312 4988 5364
rect 5040 5352 5046 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 5040 5324 5365 5352
rect 5040 5312 5046 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 5994 5312 6000 5364
rect 6052 5312 6058 5364
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 8110 5352 8116 5364
rect 8067 5324 8116 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 8846 5312 8852 5364
rect 8904 5352 8910 5364
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8904 5324 8953 5352
rect 8904 5312 8910 5324
rect 8941 5321 8953 5324
rect 8987 5321 8999 5355
rect 9858 5352 9864 5364
rect 8941 5315 8999 5321
rect 9232 5324 9864 5352
rect 9122 5284 9128 5296
rect 4856 5256 7972 5284
rect 4856 5244 4862 5256
rect 7944 5228 7972 5256
rect 8036 5256 9128 5284
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 992 5188 1593 5216
rect 992 5176 998 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 3050 5216 3056 5228
rect 2455 5188 3056 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 2240 5148 2268 5179
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 3142 5176 3148 5228
rect 3200 5176 3206 5228
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 4614 5216 4620 5228
rect 4295 5188 4620 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5074 5216 5080 5228
rect 5031 5188 5080 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 2958 5148 2964 5160
rect 2240 5120 2964 5148
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3160 5148 3188 5176
rect 4908 5148 4936 5179
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5442 5216 5448 5228
rect 5307 5188 5448 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 5905 5219 5963 5225
rect 5905 5185 5917 5219
rect 5951 5185 5963 5219
rect 5905 5179 5963 5185
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5216 6147 5219
rect 6730 5216 6736 5228
rect 6135 5188 6736 5216
rect 6135 5185 6147 5188
rect 6089 5179 6147 5185
rect 5350 5148 5356 5160
rect 3160 5120 4752 5148
rect 4908 5120 5356 5148
rect 4724 5089 4752 5120
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5920 5148 5948 5179
rect 6730 5176 6736 5188
rect 6788 5216 6794 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6788 5188 6837 5216
rect 6788 5176 6794 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 6638 5148 6644 5160
rect 5920 5120 6644 5148
rect 6638 5108 6644 5120
rect 6696 5148 6702 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6696 5120 6929 5148
rect 6696 5108 6702 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7006 5108 7012 5160
rect 7064 5108 7070 5160
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 8036 5148 8064 5256
rect 8404 5225 8432 5256
rect 9122 5244 9128 5256
rect 9180 5244 9186 5296
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 7156 5120 8064 5148
rect 7156 5108 7162 5120
rect 4709 5083 4767 5089
rect 4709 5049 4721 5083
rect 4755 5049 4767 5083
rect 4709 5043 4767 5049
rect 5166 5040 5172 5092
rect 5224 5080 5230 5092
rect 6546 5080 6552 5092
rect 5224 5052 6552 5080
rect 5224 5040 5230 5052
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 6454 4972 6460 5024
rect 6512 4972 6518 5024
rect 6564 5012 6592 5040
rect 8128 5012 8156 5179
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8588 5148 8616 5179
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 8812 5188 8861 5216
rect 8812 5176 8818 5188
rect 8849 5185 8861 5188
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5216 9091 5219
rect 9232 5216 9260 5324
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 11054 5312 11060 5364
rect 11112 5312 11118 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 13357 5355 13415 5361
rect 13357 5352 13369 5355
rect 13228 5324 13369 5352
rect 13228 5312 13234 5324
rect 13357 5321 13369 5324
rect 13403 5321 13415 5355
rect 13357 5315 13415 5321
rect 15470 5312 15476 5364
rect 15528 5312 15534 5364
rect 16114 5312 16120 5364
rect 16172 5312 16178 5364
rect 16850 5312 16856 5364
rect 16908 5312 16914 5364
rect 17218 5312 17224 5364
rect 17276 5312 17282 5364
rect 9306 5244 9312 5296
rect 9364 5284 9370 5296
rect 9585 5287 9643 5293
rect 9585 5284 9597 5287
rect 9364 5256 9597 5284
rect 9364 5244 9370 5256
rect 9585 5253 9597 5256
rect 9631 5253 9643 5287
rect 9585 5247 9643 5253
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 9732 5256 10074 5284
rect 9732 5244 9738 5256
rect 11882 5244 11888 5296
rect 11940 5244 11946 5296
rect 12618 5244 12624 5296
rect 12676 5244 12682 5296
rect 13906 5284 13912 5296
rect 13740 5256 13912 5284
rect 9079 5188 9260 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 11606 5176 11612 5228
rect 11664 5176 11670 5228
rect 13740 5225 13768 5256
rect 13906 5244 13912 5256
rect 13964 5244 13970 5296
rect 13998 5244 14004 5296
rect 14056 5244 14062 5296
rect 14090 5244 14096 5296
rect 14148 5284 14154 5296
rect 16132 5284 16160 5312
rect 14148 5256 14490 5284
rect 16040 5256 16160 5284
rect 14148 5244 14154 5256
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 15838 5176 15844 5228
rect 15896 5216 15902 5228
rect 16040 5225 16068 5256
rect 16025 5219 16083 5225
rect 16025 5216 16037 5219
rect 15896 5188 16037 5216
rect 15896 5176 15902 5188
rect 16025 5185 16037 5188
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 16114 5176 16120 5228
rect 16172 5216 16178 5228
rect 16209 5219 16267 5225
rect 16209 5216 16221 5219
rect 16172 5188 16221 5216
rect 16172 5176 16178 5188
rect 16209 5185 16221 5188
rect 16255 5185 16267 5219
rect 16209 5179 16267 5185
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16724 5188 16773 5216
rect 16724 5176 16730 5188
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 16942 5176 16948 5228
rect 17000 5176 17006 5228
rect 8260 5120 8616 5148
rect 8260 5108 8266 5120
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 8996 5120 9321 5148
rect 8996 5108 9002 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 13078 5108 13084 5160
rect 13136 5148 13142 5160
rect 16684 5148 16712 5176
rect 13136 5120 16712 5148
rect 13136 5108 13142 5120
rect 6564 4984 8156 5012
rect 8389 5015 8447 5021
rect 8389 4981 8401 5015
rect 8435 5012 8447 5015
rect 9766 5012 9772 5024
rect 8435 4984 9772 5012
rect 8435 4981 8447 4984
rect 8389 4975 8447 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 16022 4972 16028 5024
rect 16080 4972 16086 5024
rect 1104 4922 18860 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 18860 4922
rect 1104 4848 18860 4870
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 6696 4780 7389 4808
rect 6696 4768 6702 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 7377 4771 7435 4777
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 8938 4808 8944 4820
rect 7616 4780 8944 4808
rect 7616 4768 7622 4780
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10781 4811 10839 4817
rect 10781 4808 10793 4811
rect 9916 4780 10793 4808
rect 9916 4768 9922 4780
rect 10781 4777 10793 4780
rect 10827 4777 10839 4811
rect 10781 4771 10839 4777
rect 11057 4811 11115 4817
rect 11057 4777 11069 4811
rect 11103 4808 11115 4811
rect 11146 4808 11152 4820
rect 11103 4780 11152 4808
rect 11103 4777 11115 4780
rect 11057 4771 11115 4777
rect 11146 4768 11152 4780
rect 11204 4808 11210 4820
rect 11333 4811 11391 4817
rect 11333 4808 11345 4811
rect 11204 4780 11345 4808
rect 11204 4768 11210 4780
rect 11333 4777 11345 4780
rect 11379 4808 11391 4811
rect 11517 4811 11575 4817
rect 11517 4808 11529 4811
rect 11379 4780 11529 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11517 4777 11529 4780
rect 11563 4808 11575 4811
rect 11606 4808 11612 4820
rect 11563 4780 11612 4808
rect 11563 4777 11575 4780
rect 11517 4771 11575 4777
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 11701 4811 11759 4817
rect 11701 4777 11713 4811
rect 11747 4808 11759 4811
rect 12618 4808 12624 4820
rect 11747 4780 12624 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 13078 4808 13084 4820
rect 12943 4780 13084 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 4798 4700 4804 4752
rect 4856 4700 4862 4752
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 7064 4712 8156 4740
rect 7064 4700 7070 4712
rect 3326 4632 3332 4684
rect 3384 4632 3390 4684
rect 4816 4672 4844 4700
rect 4264 4644 4844 4672
rect 5905 4675 5963 4681
rect 1670 4564 1676 4616
rect 1728 4564 1734 4616
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 1946 4604 1952 4616
rect 1903 4576 1952 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 3418 4604 3424 4616
rect 3283 4576 3424 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 4264 4613 4292 4644
rect 5905 4641 5917 4675
rect 5951 4672 5963 4675
rect 6454 4672 6460 4684
rect 5951 4644 6460 4672
rect 5951 4641 5963 4644
rect 5905 4635 5963 4641
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 6914 4672 6920 4684
rect 6696 4644 6920 4672
rect 6696 4632 6702 4644
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7024 4644 8033 4672
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 5166 4604 5172 4616
rect 4847 4576 5172 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 5626 4564 5632 4616
rect 5684 4564 5690 4616
rect 7024 4590 7052 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 7926 4564 7932 4616
rect 7984 4564 7990 4616
rect 8128 4613 8156 4712
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 8720 4644 9321 4672
rect 8720 4632 8726 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 12434 4672 12440 4684
rect 9309 4635 9367 4641
rect 11716 4644 12440 4672
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8202 4604 8208 4616
rect 8159 4576 8208 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8938 4564 8944 4616
rect 8996 4604 9002 4616
rect 11716 4613 11744 4644
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 9033 4607 9091 4613
rect 9033 4604 9045 4607
rect 8996 4576 9045 4604
rect 8996 4564 9002 4576
rect 9033 4573 9045 4576
rect 9079 4573 9091 4607
rect 9033 4567 9091 4573
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 11882 4564 11888 4616
rect 11940 4564 11946 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 11992 4576 12725 4604
rect 3145 4539 3203 4545
rect 3145 4505 3157 4539
rect 3191 4536 3203 4539
rect 3602 4536 3608 4548
rect 3191 4508 3608 4536
rect 3191 4505 3203 4508
rect 3145 4499 3203 4505
rect 3602 4496 3608 4508
rect 3660 4496 3666 4548
rect 4522 4536 4528 4548
rect 4448 4508 4528 4536
rect 1854 4428 1860 4480
rect 1912 4468 1918 4480
rect 2041 4471 2099 4477
rect 2041 4468 2053 4471
rect 1912 4440 2053 4468
rect 1912 4428 1918 4440
rect 2041 4437 2053 4440
rect 2087 4437 2099 4471
rect 2041 4431 2099 4437
rect 2774 4428 2780 4480
rect 2832 4428 2838 4480
rect 4448 4477 4476 4508
rect 4522 4496 4528 4508
rect 4580 4536 4586 4548
rect 5258 4536 5264 4548
rect 4580 4508 5264 4536
rect 4580 4496 4586 4508
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4437 4491 4471
rect 4433 4431 4491 4437
rect 4706 4428 4712 4480
rect 4764 4468 4770 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 4764 4440 4997 4468
rect 4764 4428 4770 4440
rect 4985 4437 4997 4440
rect 5031 4468 5043 4471
rect 6914 4468 6920 4480
rect 5031 4440 6920 4468
rect 5031 4437 5043 4440
rect 4985 4431 5043 4437
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7558 4428 7564 4480
rect 7616 4428 7622 4480
rect 7944 4468 7972 4564
rect 9766 4496 9772 4548
rect 9824 4496 9830 4548
rect 11992 4468 12020 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 12253 4539 12311 4545
rect 12253 4505 12265 4539
rect 12299 4536 12311 4539
rect 12912 4536 12940 4771
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 13906 4808 13912 4820
rect 13679 4780 13912 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15933 4811 15991 4817
rect 15933 4808 15945 4811
rect 15252 4780 15945 4808
rect 15252 4768 15258 4780
rect 15933 4777 15945 4780
rect 15979 4777 15991 4811
rect 15933 4771 15991 4777
rect 13924 4672 13952 4768
rect 14185 4675 14243 4681
rect 14185 4672 14197 4675
rect 13924 4644 14197 4672
rect 14185 4641 14197 4644
rect 14231 4641 14243 4675
rect 14185 4635 14243 4641
rect 12299 4508 12940 4536
rect 12299 4505 12311 4508
rect 12253 4499 12311 4505
rect 14366 4496 14372 4548
rect 14424 4536 14430 4548
rect 14461 4539 14519 4545
rect 14461 4536 14473 4539
rect 14424 4508 14473 4536
rect 14424 4496 14430 4508
rect 14461 4505 14473 4508
rect 14507 4505 14519 4539
rect 16022 4536 16028 4548
rect 15686 4508 16028 4536
rect 14461 4499 14519 4505
rect 16022 4496 16028 4508
rect 16080 4496 16086 4548
rect 7944 4440 12020 4468
rect 12345 4471 12403 4477
rect 12345 4437 12357 4471
rect 12391 4468 12403 4471
rect 12434 4468 12440 4480
rect 12391 4440 12440 4468
rect 12391 4437 12403 4440
rect 12345 4431 12403 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 1104 4378 18860 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 16214 4378
rect 16266 4326 16278 4378
rect 16330 4326 16342 4378
rect 16394 4326 16406 4378
rect 16458 4326 16470 4378
rect 16522 4326 18860 4378
rect 1104 4304 18860 4326
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 4249 4267 4307 4273
rect 4249 4264 4261 4267
rect 3476 4236 4261 4264
rect 3476 4224 3482 4236
rect 4249 4233 4261 4236
rect 4295 4233 4307 4267
rect 4249 4227 4307 4233
rect 6641 4267 6699 4273
rect 6641 4233 6653 4267
rect 6687 4264 6699 4267
rect 6687 4236 7696 4264
rect 6687 4233 6699 4236
rect 6641 4227 6699 4233
rect 2774 4156 2780 4208
rect 2832 4156 2838 4208
rect 5626 4196 5632 4208
rect 4002 4168 4660 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1762 4128 1768 4140
rect 1719 4100 1768 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 1762 4088 1768 4100
rect 1820 4088 1826 4140
rect 1854 4088 1860 4140
rect 1912 4088 1918 4140
rect 2038 4088 2044 4140
rect 2096 4088 2102 4140
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2314 4128 2320 4140
rect 2179 4100 2320 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 4522 4088 4528 4140
rect 4580 4088 4586 4140
rect 4632 4137 4660 4168
rect 5276 4168 5632 4196
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 4706 4088 4712 4140
rect 4764 4088 4770 4140
rect 5276 4128 5304 4168
rect 5626 4156 5632 4168
rect 5684 4196 5690 4208
rect 6822 4196 6828 4208
rect 5684 4168 6828 4196
rect 5684 4156 5690 4168
rect 6822 4156 6828 4168
rect 6880 4196 6886 4208
rect 7558 4196 7564 4208
rect 6880 4168 7564 4196
rect 6880 4156 6886 4168
rect 4908 4100 5304 4128
rect 5353 4131 5411 4137
rect 4908 4069 4936 4100
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4128 6791 4131
rect 7006 4128 7012 4140
rect 6779 4100 7012 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 4893 4063 4951 4069
rect 4893 4060 4905 4063
rect 2547 4032 4905 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 4893 4029 4905 4032
rect 4939 4029 4951 4063
rect 4893 4023 4951 4029
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5368 3992 5396 4091
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 6362 4060 6368 4072
rect 5491 4032 6368 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 6564 4060 6592 4091
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7208 4137 7236 4168
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 7668 4196 7696 4236
rect 11146 4224 11152 4276
rect 11204 4224 11210 4276
rect 13633 4267 13691 4273
rect 13633 4233 13645 4267
rect 13679 4264 13691 4267
rect 13906 4264 13912 4276
rect 13679 4236 13912 4264
rect 13679 4233 13691 4236
rect 13633 4227 13691 4233
rect 7668 4168 7958 4196
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9640 4100 9689 4128
rect 9640 4088 9646 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 10134 4088 10140 4140
rect 10192 4088 10198 4140
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 7098 4060 7104 4072
rect 6564 4032 7104 4060
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 7466 4020 7472 4072
rect 7524 4020 7530 4072
rect 8110 4020 8116 4072
rect 8168 4060 8174 4072
rect 9214 4060 9220 4072
rect 8168 4032 9220 4060
rect 8168 4020 8174 4032
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 9456 4032 9505 4060
rect 9456 4020 9462 4032
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9493 4023 9551 4029
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 10704 4060 10732 4091
rect 9824 4032 10732 4060
rect 9824 4020 9830 4032
rect 5224 3964 5396 3992
rect 9232 3992 9260 4020
rect 10888 3992 10916 4091
rect 11808 4060 11836 4091
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 13832 4137 13860 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 15318 4168 16252 4196
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 11940 4100 11989 4128
rect 11940 4088 11946 4100
rect 11977 4097 11989 4100
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 12434 4060 12440 4072
rect 11808 4032 12440 4060
rect 12434 4020 12440 4032
rect 12492 4060 12498 4072
rect 13078 4060 13084 4072
rect 12492 4032 13084 4060
rect 12492 4020 12498 4032
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 9232 3964 10916 3992
rect 5224 3952 5230 3964
rect 11146 3952 11152 4004
rect 11204 3992 11210 4004
rect 12066 3992 12072 4004
rect 11204 3964 12072 3992
rect 11204 3952 11210 3964
rect 12066 3952 12072 3964
rect 12124 3992 12130 4004
rect 13832 3992 13860 4091
rect 15838 4088 15844 4140
rect 15896 4128 15902 4140
rect 16224 4137 16252 4168
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15896 4100 16129 4128
rect 15896 4088 15902 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4097 16267 4131
rect 16209 4091 16267 4097
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16574 4128 16580 4140
rect 16347 4100 16580 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 16574 4088 16580 4100
rect 16632 4128 16638 4140
rect 16942 4128 16948 4140
rect 16632 4100 16948 4128
rect 16632 4088 16638 4100
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17126 4088 17132 4140
rect 17184 4088 17190 4140
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 17221 4063 17279 4069
rect 14139 4032 16804 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 16776 4001 16804 4032
rect 17221 4029 17233 4063
rect 17267 4029 17279 4063
rect 17221 4023 17279 4029
rect 12124 3964 13860 3992
rect 16761 3995 16819 4001
rect 12124 3952 12130 3964
rect 16761 3961 16773 3995
rect 16807 3961 16819 3995
rect 16761 3955 16819 3961
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 3016 3896 5641 3924
rect 3016 3884 3022 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 9766 3924 9772 3936
rect 8076 3896 9772 3924
rect 8076 3884 8082 3896
rect 9766 3884 9772 3896
rect 9824 3924 9830 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9824 3896 9873 3924
rect 9824 3884 9830 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10008 3896 10333 3924
rect 10008 3884 10014 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 10778 3884 10784 3936
rect 10836 3884 10842 3936
rect 11790 3884 11796 3936
rect 11848 3884 11854 3936
rect 15565 3927 15623 3933
rect 15565 3893 15577 3927
rect 15611 3924 15623 3927
rect 16666 3924 16672 3936
rect 15611 3896 16672 3924
rect 15611 3893 15623 3896
rect 15565 3887 15623 3893
rect 16666 3884 16672 3896
rect 16724 3924 16730 3936
rect 17236 3924 17264 4023
rect 17402 4020 17408 4072
rect 17460 4020 17466 4072
rect 16724 3896 17264 3924
rect 16724 3884 16730 3896
rect 1104 3834 18860 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 18860 3834
rect 1104 3760 18860 3782
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 2866 3720 2872 3732
rect 2823 3692 2872 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5445 3723 5503 3729
rect 5445 3720 5457 3723
rect 5132 3692 5457 3720
rect 5132 3680 5138 3692
rect 5445 3689 5457 3692
rect 5491 3689 5503 3723
rect 5445 3683 5503 3689
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 7524 3692 7665 3720
rect 7524 3680 7530 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 7653 3683 7711 3689
rect 8018 3680 8024 3732
rect 8076 3680 8082 3732
rect 10134 3720 10140 3732
rect 9416 3692 10140 3720
rect 1946 3612 1952 3664
rect 2004 3652 2010 3664
rect 5169 3655 5227 3661
rect 5169 3652 5181 3655
rect 2004 3624 5181 3652
rect 2004 3612 2010 3624
rect 5169 3621 5181 3624
rect 5215 3621 5227 3655
rect 5169 3615 5227 3621
rect 5350 3612 5356 3664
rect 5408 3652 5414 3664
rect 7193 3655 7251 3661
rect 7193 3652 7205 3655
rect 5408 3624 7205 3652
rect 5408 3612 5414 3624
rect 7193 3621 7205 3624
rect 7239 3621 7251 3655
rect 9416 3652 9444 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 12161 3723 12219 3729
rect 12161 3720 12173 3723
rect 12124 3692 12173 3720
rect 12124 3680 12130 3692
rect 12161 3689 12173 3692
rect 12207 3689 12219 3723
rect 12161 3683 12219 3689
rect 13725 3723 13783 3729
rect 13725 3689 13737 3723
rect 13771 3720 13783 3723
rect 14918 3720 14924 3732
rect 13771 3692 14924 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 7193 3615 7251 3621
rect 7852 3624 9444 3652
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 2133 3587 2191 3593
rect 2133 3584 2145 3587
rect 1912 3556 2145 3584
rect 1912 3544 1918 3556
rect 2133 3553 2145 3556
rect 2179 3553 2191 3587
rect 2133 3547 2191 3553
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2501 3587 2559 3593
rect 2501 3584 2513 3587
rect 2372 3556 2513 3584
rect 2372 3544 2378 3556
rect 2501 3553 2513 3556
rect 2547 3553 2559 3587
rect 2501 3547 2559 3553
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 4764 3556 5672 3584
rect 4764 3544 4770 3556
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1670 3516 1676 3528
rect 1360 3488 1676 3516
rect 1360 3476 1366 3488
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 2096 3488 2421 3516
rect 2096 3476 2102 3488
rect 2409 3485 2421 3488
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 4798 3476 4804 3528
rect 4856 3525 4862 3528
rect 5644 3525 5672 3556
rect 4856 3519 4905 3525
rect 4856 3485 4859 3519
rect 4893 3516 4905 3519
rect 5629 3519 5687 3525
rect 4893 3488 5028 3516
rect 4893 3485 4905 3488
rect 4856 3479 4905 3485
rect 4856 3476 4862 3479
rect 2618 3451 2676 3457
rect 2618 3417 2630 3451
rect 2664 3448 2676 3451
rect 3694 3448 3700 3460
rect 2664 3420 3700 3448
rect 2664 3417 2676 3420
rect 2618 3411 2676 3417
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 5000 3448 5028 3488
rect 5629 3485 5641 3519
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 5736 3448 5764 3479
rect 5902 3476 5908 3528
rect 5960 3476 5966 3528
rect 5994 3476 6000 3528
rect 6052 3476 6058 3528
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 6979 3519 7037 3525
rect 6979 3485 6991 3519
rect 7025 3516 7037 3519
rect 7742 3516 7748 3528
rect 7025 3488 7748 3516
rect 7025 3485 7037 3488
rect 6979 3479 7037 3485
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 7852 3525 7880 3624
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 9950 3652 9956 3664
rect 9548 3624 9956 3652
rect 9548 3612 9554 3624
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 8110 3544 8116 3596
rect 8168 3544 8174 3596
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 11885 3587 11943 3593
rect 11885 3584 11897 3587
rect 9456 3556 11897 3584
rect 9456 3544 9462 3556
rect 9508 3525 9536 3556
rect 11885 3553 11897 3556
rect 11931 3553 11943 3587
rect 13740 3584 13768 3683
rect 14918 3680 14924 3692
rect 14976 3720 14982 3732
rect 16574 3720 16580 3732
rect 14976 3692 16580 3720
rect 14976 3680 14982 3692
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 17034 3680 17040 3732
rect 17092 3680 17098 3732
rect 17313 3655 17371 3661
rect 17313 3621 17325 3655
rect 17359 3621 17371 3655
rect 17313 3615 17371 3621
rect 11885 3547 11943 3553
rect 13280 3556 13768 3584
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 7837 3479 7895 3485
rect 7944 3488 9505 3516
rect 5000 3420 5764 3448
rect 1765 3383 1823 3389
rect 1765 3349 1777 3383
rect 1811 3380 1823 3383
rect 1854 3380 1860 3392
rect 1811 3352 1860 3380
rect 1811 3349 1823 3352
rect 1765 3343 1823 3349
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 7944 3380 7972 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 9582 3476 9588 3528
rect 9640 3476 9646 3528
rect 9674 3476 9680 3528
rect 9732 3476 9738 3528
rect 9861 3519 9919 3525
rect 9861 3485 9873 3519
rect 9907 3516 9919 3519
rect 9950 3516 9956 3528
rect 9907 3488 9956 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 13078 3476 13084 3528
rect 13136 3476 13142 3528
rect 13280 3525 13308 3556
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 14185 3587 14243 3593
rect 14185 3584 14197 3587
rect 13964 3556 14197 3584
rect 13964 3544 13970 3556
rect 14185 3553 14197 3556
rect 14231 3553 14243 3587
rect 14185 3547 14243 3553
rect 14461 3587 14519 3593
rect 14461 3553 14473 3587
rect 14507 3584 14519 3587
rect 17328 3584 17356 3615
rect 14507 3556 17356 3584
rect 14507 3553 14519 3556
rect 14461 3547 14519 3553
rect 17402 3544 17408 3596
rect 17460 3584 17466 3596
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17460 3556 17877 3584
rect 17460 3544 17466 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 13265 3519 13323 3525
rect 13265 3485 13277 3519
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 13556 3488 14044 3516
rect 9217 3451 9275 3457
rect 9217 3417 9229 3451
rect 9263 3448 9275 3451
rect 10413 3451 10471 3457
rect 10413 3448 10425 3451
rect 9263 3420 10425 3448
rect 9263 3417 9275 3420
rect 9217 3411 9275 3417
rect 10413 3417 10425 3420
rect 10459 3417 10471 3451
rect 11790 3448 11796 3460
rect 11638 3420 11796 3448
rect 10413 3411 10471 3417
rect 11790 3408 11796 3420
rect 11848 3408 11854 3460
rect 13173 3451 13231 3457
rect 13173 3417 13185 3451
rect 13219 3448 13231 3451
rect 13556 3448 13584 3488
rect 13219 3420 13584 3448
rect 13633 3451 13691 3457
rect 13219 3417 13231 3420
rect 13173 3411 13231 3417
rect 13633 3417 13645 3451
rect 13679 3417 13691 3451
rect 13633 3411 13691 3417
rect 6788 3352 7972 3380
rect 6788 3340 6794 3352
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13648 3380 13676 3411
rect 13044 3352 13676 3380
rect 14016 3380 14044 3488
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16393 3519 16451 3525
rect 16393 3516 16405 3519
rect 16080 3488 16405 3516
rect 16080 3476 16086 3488
rect 16393 3485 16405 3488
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 16666 3476 16672 3528
rect 16724 3516 16730 3528
rect 16761 3519 16819 3525
rect 16761 3516 16773 3519
rect 16724 3488 16773 3516
rect 16724 3476 16730 3488
rect 16761 3485 16773 3488
rect 16807 3485 16819 3519
rect 16878 3519 16936 3525
rect 16878 3516 16890 3519
rect 16761 3479 16819 3485
rect 16868 3485 16890 3516
rect 16924 3516 16936 3519
rect 17126 3516 17132 3528
rect 16924 3488 17132 3516
rect 16924 3485 16936 3488
rect 16868 3479 16936 3485
rect 16868 3448 16896 3479
rect 17126 3476 17132 3488
rect 17184 3516 17190 3528
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 17184 3488 17785 3516
rect 17184 3476 17190 3488
rect 17773 3485 17785 3488
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 17681 3451 17739 3457
rect 17681 3448 17693 3451
rect 14568 3420 14950 3448
rect 15948 3420 16896 3448
rect 16960 3420 17693 3448
rect 14568 3380 14596 3420
rect 15948 3389 15976 3420
rect 14016 3352 14596 3380
rect 15933 3383 15991 3389
rect 13044 3340 13050 3352
rect 15933 3349 15945 3383
rect 15979 3349 15991 3383
rect 15933 3343 15991 3349
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 16960 3380 16988 3420
rect 17681 3417 17693 3420
rect 17727 3417 17739 3451
rect 17681 3411 17739 3417
rect 16724 3352 16988 3380
rect 16724 3340 16730 3352
rect 1104 3290 18860 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 16214 3290
rect 16266 3238 16278 3290
rect 16330 3238 16342 3290
rect 16394 3238 16406 3290
rect 16458 3238 16470 3290
rect 16522 3238 18860 3290
rect 1104 3216 18860 3238
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 2593 3179 2651 3185
rect 2593 3176 2605 3179
rect 2372 3148 2605 3176
rect 2372 3136 2378 3148
rect 2593 3145 2605 3148
rect 2639 3145 2651 3179
rect 2593 3139 2651 3145
rect 3694 3136 3700 3188
rect 3752 3136 3758 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 4764 3148 5580 3176
rect 4764 3136 4770 3148
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 4798 3108 4804 3120
rect 1811 3080 2360 3108
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2130 3040 2136 3052
rect 1719 3012 2136 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 2332 3049 2360 3080
rect 3436 3080 4804 3108
rect 3436 3052 3464 3080
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 5552 3117 5580 3148
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 5960 3148 7021 3176
rect 5960 3136 5966 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 7009 3139 7067 3145
rect 7742 3136 7748 3188
rect 7800 3176 7806 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 7800 3148 8033 3176
rect 7800 3136 7806 3148
rect 8021 3145 8033 3148
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 8849 3179 8907 3185
rect 8849 3145 8861 3179
rect 8895 3176 8907 3179
rect 9030 3176 9036 3188
rect 8895 3148 9036 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 9030 3136 9036 3148
rect 9088 3176 9094 3188
rect 9582 3176 9588 3188
rect 9088 3148 9588 3176
rect 9088 3136 9094 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 9732 3148 9873 3176
rect 9732 3136 9738 3148
rect 9861 3145 9873 3148
rect 9907 3145 9919 3179
rect 9861 3139 9919 3145
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 13449 3179 13507 3185
rect 13449 3176 13461 3179
rect 11011 3148 13461 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 13449 3145 13461 3148
rect 13495 3145 13507 3179
rect 13449 3139 13507 3145
rect 13725 3179 13783 3185
rect 13725 3145 13737 3179
rect 13771 3176 13783 3179
rect 13906 3176 13912 3188
rect 13771 3148 13912 3176
rect 13771 3145 13783 3148
rect 13725 3139 13783 3145
rect 5537 3111 5595 3117
rect 5537 3077 5549 3111
rect 5583 3077 5595 3111
rect 6730 3108 6736 3120
rect 5537 3071 5595 3077
rect 6656 3080 6736 3108
rect 5448 3052 5500 3058
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2774 3040 2780 3052
rect 2455 3012 2780 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 2240 2972 2268 3003
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3418 3000 3424 3052
rect 3476 3000 3482 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4614 3040 4620 3052
rect 4387 3012 4620 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 1360 2944 3709 2972
rect 1360 2932 1366 2944
rect 3697 2941 3709 2944
rect 3743 2941 3755 2975
rect 3697 2935 3755 2941
rect 4172 2904 4200 3003
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 6656 3049 6684 3080
rect 6730 3068 6736 3080
rect 6788 3108 6794 3120
rect 7834 3108 7840 3120
rect 6788 3080 7840 3108
rect 6788 3068 6794 3080
rect 7668 3049 7696 3080
rect 7834 3068 7840 3080
rect 7892 3108 7898 3120
rect 8478 3108 8484 3120
rect 7892 3080 8484 3108
rect 7892 3068 7898 3080
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 8662 3068 8668 3120
rect 8720 3117 8726 3120
rect 8720 3111 8739 3117
rect 8727 3077 8739 3111
rect 10980 3108 11008 3139
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 15657 3179 15715 3185
rect 15657 3145 15669 3179
rect 15703 3176 15715 3179
rect 16666 3176 16672 3188
rect 15703 3148 16672 3176
rect 15703 3145 15715 3148
rect 15657 3139 15715 3145
rect 16666 3136 16672 3148
rect 16724 3176 16730 3188
rect 16724 3148 16988 3176
rect 16724 3136 16730 3148
rect 12066 3108 12072 3120
rect 8720 3071 8739 3077
rect 8772 3080 11008 3108
rect 11716 3080 12072 3108
rect 8720 3068 8726 3071
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3040 6883 3043
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 6871 3012 7481 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 5448 2994 5500 3000
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 5074 2972 5080 2984
rect 5031 2944 5080 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 7484 2972 7512 3003
rect 7944 2972 7972 3003
rect 8772 2972 8800 3080
rect 11716 3052 11744 3080
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 12986 3068 12992 3120
rect 13044 3068 13050 3120
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 9272 3012 9505 3040
rect 9272 3000 9278 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9647 3043 9705 3049
rect 9647 3009 9659 3043
rect 9693 3040 9705 3043
rect 9766 3040 9772 3052
rect 9693 3012 9772 3040
rect 9693 3009 9705 3012
rect 9647 3003 9705 3009
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 9876 3012 10885 3040
rect 9876 2972 9904 3012
rect 10873 3009 10885 3012
rect 10919 3040 10931 3043
rect 11238 3040 11244 3052
rect 10919 3012 11244 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 13924 3049 13952 3136
rect 16301 3111 16359 3117
rect 16301 3108 16313 3111
rect 15410 3080 16313 3108
rect 16301 3077 16313 3080
rect 16347 3077 16359 3111
rect 16301 3071 16359 3077
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 15838 3040 15844 3052
rect 15620 3012 15844 3040
rect 15620 3000 15626 3012
rect 15838 3000 15844 3012
rect 15896 3040 15902 3052
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 15896 3012 16221 3040
rect 15896 3000 15902 3012
rect 16209 3009 16221 3012
rect 16255 3009 16267 3043
rect 16209 3003 16267 3009
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3040 16451 3043
rect 16574 3040 16580 3052
rect 16439 3012 16580 3040
rect 16439 3009 16451 3012
rect 16393 3003 16451 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 16960 3049 16988 3148
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 17099 3043 17157 3049
rect 17099 3009 17111 3043
rect 17145 3040 17157 3043
rect 17402 3040 17408 3052
rect 17145 3012 17408 3040
rect 17145 3009 17157 3012
rect 17099 3003 17157 3009
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 17678 3000 17684 3052
rect 17736 3000 17742 3052
rect 7484 2944 8800 2972
rect 9646 2944 9904 2972
rect 4172 2876 5304 2904
rect 5276 2848 5304 2876
rect 8478 2864 8484 2916
rect 8536 2904 8542 2916
rect 9646 2904 9674 2944
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 10284 2944 11069 2972
rect 10284 2932 10290 2944
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 8536 2876 9674 2904
rect 10505 2907 10563 2913
rect 8536 2864 8542 2876
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 10962 2904 10968 2916
rect 10551 2876 10968 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 2130 2796 2136 2848
rect 2188 2836 2194 2848
rect 3513 2839 3571 2845
rect 3513 2836 3525 2839
rect 2188 2808 3525 2836
rect 2188 2796 2194 2808
rect 3513 2805 3525 2808
rect 3559 2805 3571 2839
rect 3513 2799 3571 2805
rect 3970 2796 3976 2848
rect 4028 2836 4034 2848
rect 4157 2839 4215 2845
rect 4157 2836 4169 2839
rect 4028 2808 4169 2836
rect 4028 2796 4034 2808
rect 4157 2805 4169 2808
rect 4203 2805 4215 2839
rect 4157 2799 4215 2805
rect 5258 2796 5264 2848
rect 5316 2836 5322 2848
rect 7006 2836 7012 2848
rect 5316 2808 7012 2836
rect 5316 2796 5322 2808
rect 7006 2796 7012 2808
rect 7064 2836 7070 2848
rect 7190 2836 7196 2848
rect 7064 2808 7196 2836
rect 7064 2796 7070 2808
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 7466 2796 7472 2848
rect 7524 2796 7530 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8352 2808 8677 2836
rect 8352 2796 8358 2808
rect 8665 2805 8677 2808
rect 8711 2836 8723 2839
rect 8754 2836 8760 2848
rect 8711 2808 8760 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 11072 2836 11100 2935
rect 11146 2932 11152 2984
rect 11204 2972 11210 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11204 2944 11989 2972
rect 11204 2932 11210 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 14185 2975 14243 2981
rect 12124 2944 14044 2972
rect 12124 2932 12130 2944
rect 12066 2836 12072 2848
rect 11072 2808 12072 2836
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 14016 2836 14044 2944
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 14231 2944 17325 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 16022 2836 16028 2848
rect 14016 2808 16028 2836
rect 16022 2796 16028 2808
rect 16080 2836 16086 2848
rect 17420 2836 17448 3000
rect 17773 2839 17831 2845
rect 17773 2836 17785 2839
rect 16080 2808 17785 2836
rect 16080 2796 16086 2808
rect 17773 2805 17785 2808
rect 17819 2805 17831 2839
rect 17773 2799 17831 2805
rect 1104 2746 18860 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 18860 2746
rect 1104 2672 18860 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2038 2632 2044 2644
rect 1995 2604 2044 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2593 2635 2651 2641
rect 2593 2632 2605 2635
rect 2188 2604 2605 2632
rect 2188 2592 2194 2604
rect 2593 2601 2605 2604
rect 2639 2601 2651 2635
rect 2593 2595 2651 2601
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 2832 2604 3985 2632
rect 2832 2592 2838 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 5166 2632 5172 2644
rect 4571 2604 5172 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 5994 2632 6000 2644
rect 5859 2604 6000 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 3418 2524 3424 2576
rect 3476 2524 3482 2576
rect 1946 2496 1952 2508
rect 1780 2468 1952 2496
rect 1780 2437 1808 2468
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 5828 2496 5856 2595
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6362 2592 6368 2644
rect 6420 2592 6426 2644
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 9858 2632 9864 2644
rect 6972 2604 9864 2632
rect 6972 2592 6978 2604
rect 7837 2567 7895 2573
rect 2608 2468 3280 2496
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 1854 2388 1860 2440
rect 1912 2428 1918 2440
rect 2608 2437 2636 2468
rect 2593 2431 2651 2437
rect 1912 2400 1957 2428
rect 1912 2388 1918 2400
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 2958 2428 2964 2440
rect 2823 2400 2964 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 2958 2388 2964 2400
rect 3016 2428 3022 2440
rect 3252 2437 3280 2468
rect 4540 2468 5856 2496
rect 6472 2536 7788 2564
rect 3145 2431 3203 2437
rect 3145 2428 3157 2431
rect 3016 2400 3157 2428
rect 3016 2388 3022 2400
rect 3145 2397 3157 2400
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3694 2428 3700 2440
rect 3283 2400 3700 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3160 2360 3188 2391
rect 3694 2388 3700 2400
rect 3752 2428 3758 2440
rect 3881 2431 3939 2437
rect 3881 2428 3893 2431
rect 3752 2400 3893 2428
rect 3752 2388 3758 2400
rect 3881 2397 3893 2400
rect 3927 2397 3939 2431
rect 3881 2391 3939 2397
rect 4062 2388 4068 2440
rect 4120 2388 4126 2440
rect 4540 2437 4568 2468
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4764 2400 4813 2428
rect 4764 2388 4770 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5074 2388 5080 2440
rect 5132 2428 5138 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5132 2400 5457 2428
rect 5132 2388 5138 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 4080 2360 4108 2388
rect 3160 2332 4108 2360
rect 5460 2360 5488 2391
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 5592 2400 5641 2428
rect 5592 2388 5598 2400
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 5902 2388 5908 2440
rect 5960 2428 5966 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5960 2400 6377 2428
rect 5960 2388 5966 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 6472 2360 6500 2536
rect 7466 2496 7472 2508
rect 6564 2468 7472 2496
rect 6564 2437 6592 2468
rect 7466 2456 7472 2468
rect 7524 2456 7530 2508
rect 7760 2496 7788 2536
rect 7837 2533 7849 2567
rect 7883 2564 7895 2567
rect 9125 2567 9183 2573
rect 9125 2564 9137 2567
rect 7883 2536 9137 2564
rect 7883 2533 7895 2536
rect 7837 2527 7895 2533
rect 9125 2533 9137 2536
rect 9171 2533 9183 2567
rect 9125 2527 9183 2533
rect 8018 2496 8024 2508
rect 7760 2468 8024 2496
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 9324 2505 9352 2604
rect 9858 2592 9864 2604
rect 9916 2632 9922 2644
rect 10778 2632 10784 2644
rect 9916 2604 10784 2632
rect 9916 2592 9922 2604
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11296 2604 11621 2632
rect 11296 2592 11302 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 12986 2592 12992 2644
rect 13044 2592 13050 2644
rect 16025 2567 16083 2573
rect 16025 2564 16037 2567
rect 14200 2536 16037 2564
rect 9309 2499 9367 2505
rect 9309 2465 9321 2499
rect 9355 2465 9367 2499
rect 10134 2496 10140 2508
rect 9309 2459 9367 2465
rect 9876 2468 10140 2496
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7006 2428 7012 2440
rect 6963 2400 7012 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7616 2400 8125 2428
rect 7616 2388 7622 2400
rect 8113 2397 8125 2400
rect 8159 2428 8171 2431
rect 8662 2428 8668 2440
rect 8159 2400 8668 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9030 2388 9036 2440
rect 9088 2388 9094 2440
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9876 2437 9904 2468
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10226 2456 10232 2508
rect 10284 2496 10290 2508
rect 14200 2496 14228 2536
rect 16025 2533 16037 2536
rect 16071 2564 16083 2567
rect 17678 2564 17684 2576
rect 16071 2536 17684 2564
rect 16071 2533 16083 2536
rect 16025 2527 16083 2533
rect 17678 2524 17684 2536
rect 17736 2524 17742 2576
rect 15562 2496 15568 2508
rect 10284 2468 14228 2496
rect 14292 2468 15568 2496
rect 10284 2456 10290 2468
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9732 2400 9873 2428
rect 9732 2388 9738 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 12986 2388 12992 2440
rect 13044 2388 13050 2440
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 14185 2431 14243 2437
rect 14185 2397 14197 2431
rect 14231 2428 14243 2431
rect 14292 2428 14320 2468
rect 14384 2437 14504 2438
rect 14844 2437 14872 2468
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 15746 2456 15752 2508
rect 15804 2456 15810 2508
rect 14231 2400 14320 2428
rect 14369 2431 14504 2437
rect 14231 2397 14243 2400
rect 14185 2391 14243 2397
rect 14369 2397 14381 2431
rect 14415 2410 14504 2431
rect 14415 2397 14427 2410
rect 14369 2391 14427 2397
rect 5460 2332 6500 2360
rect 7834 2320 7840 2372
rect 7892 2320 7898 2372
rect 8018 2320 8024 2372
rect 8076 2360 8082 2372
rect 8294 2360 8300 2372
rect 8076 2332 8300 2360
rect 8076 2320 8082 2332
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 8481 2363 8539 2369
rect 8481 2329 8493 2363
rect 8527 2329 8539 2363
rect 8481 2323 8539 2329
rect 4709 2295 4767 2301
rect 4709 2261 4721 2295
rect 4755 2292 4767 2295
rect 4798 2292 4804 2304
rect 4755 2264 4804 2292
rect 4755 2261 4767 2264
rect 4709 2255 4767 2261
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 6546 2252 6552 2304
rect 6604 2292 6610 2304
rect 6914 2292 6920 2304
rect 6604 2264 6920 2292
rect 6604 2252 6610 2264
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7006 2252 7012 2304
rect 7064 2252 7070 2304
rect 7466 2252 7472 2304
rect 7524 2292 7530 2304
rect 8110 2292 8116 2304
rect 7524 2264 8116 2292
rect 7524 2252 7530 2264
rect 8110 2252 8116 2264
rect 8168 2292 8174 2304
rect 8496 2292 8524 2323
rect 10134 2320 10140 2372
rect 10192 2320 10198 2372
rect 10870 2320 10876 2372
rect 10928 2320 10934 2372
rect 13188 2360 13216 2391
rect 14476 2360 14504 2410
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14976 2400 15025 2428
rect 14976 2388 14982 2400
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 15528 2400 15669 2428
rect 15528 2388 15534 2400
rect 15657 2397 15669 2400
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 14936 2360 14964 2388
rect 13188 2332 14964 2360
rect 8168 2264 8524 2292
rect 9309 2295 9367 2301
rect 8168 2252 8174 2264
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 9582 2292 9588 2304
rect 9355 2264 9588 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 11698 2252 11704 2304
rect 11756 2292 11762 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11756 2264 11805 2292
rect 11756 2252 11762 2264
rect 11793 2261 11805 2264
rect 11839 2292 11851 2295
rect 11977 2295 12035 2301
rect 11977 2292 11989 2295
rect 11839 2264 11989 2292
rect 11839 2261 11851 2264
rect 11793 2255 11851 2261
rect 11977 2261 11989 2264
rect 12023 2261 12035 2295
rect 11977 2255 12035 2261
rect 13722 2252 13728 2304
rect 13780 2252 13786 2304
rect 14274 2252 14280 2304
rect 14332 2252 14338 2304
rect 14918 2252 14924 2304
rect 14976 2252 14982 2304
rect 1104 2202 18860 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 16214 2202
rect 16266 2150 16278 2202
rect 16330 2150 16342 2202
rect 16394 2150 16406 2202
rect 16458 2150 16470 2202
rect 16522 2150 18860 2202
rect 1104 2128 18860 2150
rect 3694 2048 3700 2100
rect 3752 2048 3758 2100
rect 6089 2091 6147 2097
rect 6089 2088 6101 2091
rect 4080 2060 6101 2088
rect 3970 2020 3976 2032
rect 3450 1992 3976 2020
rect 3970 1980 3976 1992
rect 4028 1980 4034 2032
rect 1946 1912 1952 1964
rect 2004 1912 2010 1964
rect 3878 1912 3884 1964
rect 3936 1952 3942 1964
rect 4080 1961 4108 2060
rect 6089 2057 6101 2060
rect 6135 2088 6147 2091
rect 6730 2088 6736 2100
rect 6135 2060 6736 2088
rect 6135 2057 6147 2060
rect 6089 2051 6147 2057
rect 6730 2048 6736 2060
rect 6788 2088 6794 2100
rect 9674 2088 9680 2100
rect 6788 2060 6914 2088
rect 6788 2048 6794 2060
rect 4798 1980 4804 2032
rect 4856 1980 4862 2032
rect 6457 2023 6515 2029
rect 6457 1989 6469 2023
rect 6503 2020 6515 2023
rect 6546 2020 6552 2032
rect 6503 1992 6552 2020
rect 6503 1989 6515 1992
rect 6457 1983 6515 1989
rect 6546 1980 6552 1992
rect 6604 1980 6610 2032
rect 6886 2020 6914 2060
rect 8404 2060 9680 2088
rect 8404 2020 8432 2060
rect 9674 2048 9680 2060
rect 9732 2048 9738 2100
rect 10870 2048 10876 2100
rect 10928 2048 10934 2100
rect 13449 2091 13507 2097
rect 13449 2057 13461 2091
rect 13495 2088 13507 2091
rect 13495 2060 14044 2088
rect 13495 2057 13507 2060
rect 13449 2051 13507 2057
rect 10594 2020 10600 2032
rect 6886 1992 8432 2020
rect 9890 1992 10600 2020
rect 8404 1964 8432 1992
rect 10594 1980 10600 1992
rect 10652 1980 10658 2032
rect 11882 1980 11888 2032
rect 11940 2020 11946 2032
rect 14016 2029 14044 2060
rect 14001 2023 14059 2029
rect 11940 1992 12466 2020
rect 11940 1980 11946 1992
rect 14001 1989 14013 2023
rect 14047 1989 14059 2023
rect 14001 1983 14059 1989
rect 14274 1980 14280 2032
rect 14332 2020 14338 2032
rect 14332 1992 14490 2020
rect 14332 1980 14338 1992
rect 4065 1955 4123 1961
rect 4065 1952 4077 1955
rect 3936 1924 4077 1952
rect 3936 1912 3942 1924
rect 4065 1921 4077 1924
rect 4111 1921 4123 1955
rect 4065 1915 4123 1921
rect 6362 1912 6368 1964
rect 6420 1952 6426 1964
rect 6638 1952 6644 1964
rect 6420 1924 6644 1952
rect 6420 1912 6426 1924
rect 6638 1912 6644 1924
rect 6696 1912 6702 1964
rect 6733 1955 6791 1961
rect 6733 1921 6745 1955
rect 6779 1952 6791 1955
rect 7466 1952 7472 1964
rect 6779 1924 7472 1952
rect 6779 1921 6791 1924
rect 6733 1915 6791 1921
rect 7466 1912 7472 1924
rect 7524 1912 7530 1964
rect 7653 1955 7711 1961
rect 7653 1921 7665 1955
rect 7699 1952 7711 1955
rect 8018 1952 8024 1964
rect 7699 1924 8024 1952
rect 7699 1921 7711 1924
rect 7653 1915 7711 1921
rect 8018 1912 8024 1924
rect 8076 1912 8082 1964
rect 8386 1912 8392 1964
rect 8444 1912 8450 1964
rect 10778 1912 10784 1964
rect 10836 1912 10842 1964
rect 10965 1955 11023 1961
rect 10965 1921 10977 1955
rect 11011 1952 11023 1955
rect 11146 1952 11152 1964
rect 11011 1924 11152 1952
rect 11011 1921 11023 1924
rect 10965 1915 11023 1921
rect 11146 1912 11152 1924
rect 11204 1952 11210 1964
rect 11606 1952 11612 1964
rect 11204 1924 11612 1952
rect 11204 1912 11210 1924
rect 11606 1912 11612 1924
rect 11664 1912 11670 1964
rect 2225 1887 2283 1893
rect 2225 1853 2237 1887
rect 2271 1884 2283 1887
rect 2590 1884 2596 1896
rect 2271 1856 2596 1884
rect 2271 1853 2283 1856
rect 2225 1847 2283 1853
rect 2590 1844 2596 1856
rect 2648 1844 2654 1896
rect 4341 1887 4399 1893
rect 4341 1853 4353 1887
rect 4387 1884 4399 1887
rect 4890 1884 4896 1896
rect 4387 1856 4896 1884
rect 4387 1853 4399 1856
rect 4341 1847 4399 1853
rect 4890 1844 4896 1856
rect 4948 1844 4954 1896
rect 7558 1884 7564 1896
rect 5368 1856 7564 1884
rect 4062 1708 4068 1760
rect 4120 1748 4126 1760
rect 5368 1748 5396 1856
rect 7558 1844 7564 1856
rect 7616 1844 7622 1896
rect 8662 1844 8668 1896
rect 8720 1844 8726 1896
rect 8754 1844 8760 1896
rect 8812 1884 8818 1896
rect 10413 1887 10471 1893
rect 10413 1884 10425 1887
rect 8812 1856 10425 1884
rect 8812 1844 8818 1856
rect 10413 1853 10425 1856
rect 10459 1853 10471 1887
rect 11698 1884 11704 1896
rect 10413 1847 10471 1853
rect 11256 1856 11704 1884
rect 5442 1776 5448 1828
rect 5500 1816 5506 1828
rect 5813 1819 5871 1825
rect 5813 1816 5825 1819
rect 5500 1788 5825 1816
rect 5500 1776 5506 1788
rect 5813 1785 5825 1788
rect 5859 1785 5871 1819
rect 5813 1779 5871 1785
rect 11256 1760 11284 1856
rect 11698 1844 11704 1856
rect 11756 1844 11762 1896
rect 11977 1887 12035 1893
rect 11977 1853 11989 1887
rect 12023 1884 12035 1887
rect 12023 1856 13676 1884
rect 12023 1853 12035 1856
rect 11977 1847 12035 1853
rect 4120 1720 5396 1748
rect 4120 1708 4126 1720
rect 6546 1708 6552 1760
rect 6604 1708 6610 1760
rect 7929 1751 7987 1757
rect 7929 1717 7941 1751
rect 7975 1748 7987 1751
rect 9766 1748 9772 1760
rect 7975 1720 9772 1748
rect 7975 1717 7987 1720
rect 7929 1711 7987 1717
rect 9766 1708 9772 1720
rect 9824 1708 9830 1760
rect 11238 1708 11244 1760
rect 11296 1708 11302 1760
rect 13648 1748 13676 1856
rect 13722 1844 13728 1896
rect 13780 1844 13786 1896
rect 14550 1748 14556 1760
rect 13648 1720 14556 1748
rect 14550 1708 14556 1720
rect 14608 1708 14614 1760
rect 15470 1708 15476 1760
rect 15528 1708 15534 1760
rect 1104 1658 18860 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 18860 1658
rect 1104 1584 18860 1606
rect 1946 1504 1952 1556
rect 2004 1544 2010 1556
rect 2317 1547 2375 1553
rect 2317 1544 2329 1547
rect 2004 1516 2329 1544
rect 2004 1504 2010 1516
rect 2317 1513 2329 1516
rect 2363 1544 2375 1547
rect 3878 1544 3884 1556
rect 2363 1516 3884 1544
rect 2363 1513 2375 1516
rect 2317 1507 2375 1513
rect 3878 1504 3884 1516
rect 3936 1504 3942 1556
rect 4249 1547 4307 1553
rect 4249 1513 4261 1547
rect 4295 1544 4307 1547
rect 4798 1544 4804 1556
rect 4295 1516 4804 1544
rect 4295 1513 4307 1516
rect 4249 1507 4307 1513
rect 4798 1504 4804 1516
rect 4856 1504 4862 1556
rect 4890 1504 4896 1556
rect 4948 1504 4954 1556
rect 6546 1504 6552 1556
rect 6604 1544 6610 1556
rect 6714 1547 6772 1553
rect 6714 1544 6726 1547
rect 6604 1516 6726 1544
rect 6604 1504 6610 1516
rect 6714 1513 6726 1516
rect 6760 1513 6772 1547
rect 6714 1507 6772 1513
rect 8110 1504 8116 1556
rect 8168 1544 8174 1556
rect 8205 1547 8263 1553
rect 8205 1544 8217 1547
rect 8168 1516 8217 1544
rect 8168 1504 8174 1516
rect 8205 1513 8217 1516
rect 8251 1513 8263 1547
rect 8205 1507 8263 1513
rect 8386 1504 8392 1556
rect 8444 1504 8450 1556
rect 8662 1504 8668 1556
rect 8720 1544 8726 1556
rect 9493 1547 9551 1553
rect 9493 1544 9505 1547
rect 8720 1516 9505 1544
rect 8720 1504 8726 1516
rect 9493 1513 9505 1516
rect 9539 1513 9551 1547
rect 9493 1507 9551 1513
rect 9674 1504 9680 1556
rect 9732 1544 9738 1556
rect 10689 1547 10747 1553
rect 10689 1544 10701 1547
rect 9732 1516 10701 1544
rect 9732 1504 9738 1516
rect 10689 1513 10701 1516
rect 10735 1544 10747 1547
rect 11238 1544 11244 1556
rect 10735 1516 11244 1544
rect 10735 1513 10747 1516
rect 10689 1507 10747 1513
rect 11238 1504 11244 1516
rect 11296 1544 11302 1556
rect 13541 1547 13599 1553
rect 13541 1544 13553 1547
rect 11296 1516 13553 1544
rect 11296 1504 11302 1516
rect 13541 1513 13553 1516
rect 13587 1544 13599 1547
rect 13722 1544 13728 1556
rect 13587 1516 13728 1544
rect 13587 1513 13599 1516
rect 13541 1507 13599 1513
rect 13722 1504 13728 1516
rect 13780 1544 13786 1556
rect 13817 1547 13875 1553
rect 13817 1544 13829 1547
rect 13780 1516 13829 1544
rect 13780 1504 13786 1516
rect 13817 1513 13829 1516
rect 13863 1513 13875 1547
rect 13817 1507 13875 1513
rect 2590 1436 2596 1488
rect 2648 1436 2654 1488
rect 10134 1436 10140 1488
rect 10192 1476 10198 1488
rect 10505 1479 10563 1485
rect 10505 1476 10517 1479
rect 10192 1448 10517 1476
rect 10192 1436 10198 1448
rect 10505 1445 10517 1448
rect 10551 1445 10563 1479
rect 10505 1439 10563 1445
rect 10594 1436 10600 1488
rect 10652 1476 10658 1488
rect 10965 1479 11023 1485
rect 10965 1476 10977 1479
rect 10652 1448 10977 1476
rect 10652 1436 10658 1448
rect 10965 1445 10977 1448
rect 11011 1445 11023 1479
rect 10965 1439 11023 1445
rect 11882 1436 11888 1488
rect 11940 1436 11946 1488
rect 3237 1411 3295 1417
rect 3237 1377 3249 1411
rect 3283 1408 3295 1411
rect 3326 1408 3332 1420
rect 3283 1380 3332 1408
rect 3283 1377 3295 1380
rect 3237 1371 3295 1377
rect 3326 1368 3332 1380
rect 3384 1408 3390 1420
rect 5445 1411 5503 1417
rect 5445 1408 5457 1411
rect 3384 1380 5457 1408
rect 3384 1368 3390 1380
rect 5445 1377 5457 1380
rect 5491 1408 5503 1411
rect 6362 1408 6368 1420
rect 5491 1380 6368 1408
rect 5491 1377 5503 1380
rect 5445 1371 5503 1377
rect 6362 1368 6368 1380
rect 6420 1368 6426 1420
rect 6457 1411 6515 1417
rect 6457 1377 6469 1411
rect 6503 1408 6515 1411
rect 6730 1408 6736 1420
rect 6503 1380 6736 1408
rect 6503 1377 6515 1380
rect 6457 1371 6515 1377
rect 6730 1368 6736 1380
rect 6788 1368 6794 1420
rect 13832 1408 13860 1507
rect 15746 1504 15752 1556
rect 15804 1544 15810 1556
rect 15933 1547 15991 1553
rect 15933 1544 15945 1547
rect 15804 1516 15945 1544
rect 15804 1504 15810 1516
rect 15933 1513 15945 1516
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 14185 1411 14243 1417
rect 14185 1408 14197 1411
rect 11164 1380 12112 1408
rect 13832 1380 14197 1408
rect 11164 1352 11192 1380
rect 1765 1343 1823 1349
rect 1765 1309 1777 1343
rect 1811 1340 1823 1343
rect 1946 1340 1952 1352
rect 1811 1312 1952 1340
rect 1811 1309 1823 1312
rect 1765 1303 1823 1309
rect 1946 1300 1952 1312
rect 2004 1300 2010 1352
rect 2958 1300 2964 1352
rect 3016 1300 3022 1352
rect 3053 1343 3111 1349
rect 3053 1309 3065 1343
rect 3099 1340 3111 1343
rect 3694 1340 3700 1352
rect 3099 1312 3700 1340
rect 3099 1309 3111 1312
rect 3053 1303 3111 1309
rect 3694 1300 3700 1312
rect 3752 1300 3758 1352
rect 4249 1343 4307 1349
rect 4249 1309 4261 1343
rect 4295 1309 4307 1343
rect 4249 1303 4307 1309
rect 4433 1343 4491 1349
rect 4433 1309 4445 1343
rect 4479 1340 4491 1343
rect 4614 1340 4620 1352
rect 4479 1312 4620 1340
rect 4479 1309 4491 1312
rect 4433 1303 4491 1309
rect 4264 1272 4292 1303
rect 4614 1300 4620 1312
rect 4672 1300 4678 1352
rect 5074 1300 5080 1352
rect 5132 1340 5138 1352
rect 5261 1343 5319 1349
rect 5261 1340 5273 1343
rect 5132 1312 5273 1340
rect 5132 1300 5138 1312
rect 5261 1309 5273 1312
rect 5307 1309 5319 1343
rect 5261 1303 5319 1309
rect 9309 1343 9367 1349
rect 9309 1309 9321 1343
rect 9355 1340 9367 1343
rect 9490 1340 9496 1352
rect 9355 1312 9496 1340
rect 9355 1309 9367 1312
rect 9309 1303 9367 1309
rect 5166 1272 5172 1284
rect 4264 1244 5172 1272
rect 5166 1232 5172 1244
rect 5224 1232 5230 1284
rect 5353 1275 5411 1281
rect 5353 1241 5365 1275
rect 5399 1272 5411 1275
rect 5442 1272 5448 1284
rect 5399 1244 5448 1272
rect 5399 1241 5411 1244
rect 5353 1235 5411 1241
rect 5442 1232 5448 1244
rect 5500 1232 5506 1284
rect 7006 1232 7012 1284
rect 7064 1272 7070 1284
rect 7064 1244 7222 1272
rect 7064 1232 7070 1244
rect 1026 1164 1032 1216
rect 1084 1204 1090 1216
rect 1949 1207 2007 1213
rect 1949 1204 1961 1207
rect 1084 1176 1961 1204
rect 1084 1164 1090 1176
rect 1949 1173 1961 1176
rect 1995 1173 2007 1207
rect 1949 1167 2007 1173
rect 6362 1164 6368 1216
rect 6420 1204 6426 1216
rect 9324 1204 9352 1303
rect 9490 1300 9496 1312
rect 9548 1300 9554 1352
rect 9766 1300 9772 1352
rect 9824 1300 9830 1352
rect 10226 1300 10232 1352
rect 10284 1300 10290 1352
rect 10321 1343 10379 1349
rect 10321 1309 10333 1343
rect 10367 1309 10379 1343
rect 10321 1303 10379 1309
rect 9582 1232 9588 1284
rect 9640 1272 9646 1284
rect 10336 1272 10364 1303
rect 10778 1300 10784 1352
rect 10836 1340 10842 1352
rect 10965 1343 11023 1349
rect 10965 1340 10977 1343
rect 10836 1312 10977 1340
rect 10836 1300 10842 1312
rect 10965 1309 10977 1312
rect 11011 1309 11023 1343
rect 10965 1303 11023 1309
rect 9640 1244 10364 1272
rect 10980 1272 11008 1303
rect 11146 1300 11152 1352
rect 11204 1300 11210 1352
rect 12084 1349 12112 1380
rect 14185 1377 14197 1380
rect 14231 1377 14243 1411
rect 14185 1371 14243 1377
rect 14461 1411 14519 1417
rect 14461 1377 14473 1411
rect 14507 1408 14519 1411
rect 15470 1408 15476 1420
rect 14507 1380 15476 1408
rect 14507 1377 14519 1380
rect 14461 1371 14519 1377
rect 15470 1368 15476 1380
rect 15528 1368 15534 1420
rect 11885 1343 11943 1349
rect 11885 1309 11897 1343
rect 11931 1309 11943 1343
rect 11885 1303 11943 1309
rect 12069 1343 12127 1349
rect 12069 1309 12081 1343
rect 12115 1309 12127 1343
rect 12069 1303 12127 1309
rect 11900 1272 11928 1303
rect 12986 1272 12992 1284
rect 10980 1244 12992 1272
rect 9640 1232 9646 1244
rect 12986 1232 12992 1244
rect 13044 1232 13050 1284
rect 14918 1232 14924 1284
rect 14976 1232 14982 1284
rect 6420 1176 9352 1204
rect 9677 1207 9735 1213
rect 6420 1164 6426 1176
rect 9677 1173 9689 1207
rect 9723 1204 9735 1207
rect 9858 1204 9864 1216
rect 9723 1176 9864 1204
rect 9723 1173 9735 1176
rect 9677 1167 9735 1173
rect 9858 1164 9864 1176
rect 9916 1164 9922 1216
rect 1104 1114 18860 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 16214 1114
rect 16266 1062 16278 1114
rect 16330 1062 16342 1114
rect 16394 1062 16406 1114
rect 16458 1062 16470 1114
rect 16522 1062 18860 1114
rect 1104 1040 18860 1062
<< via1 >>
rect 1400 14288 1452 14340
rect 7104 14288 7156 14340
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 3056 13336 3108 13388
rect 12256 13472 12308 13524
rect 6920 13336 6972 13388
rect 7840 13336 7892 13388
rect 4068 13268 4120 13320
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 4804 13132 4856 13184
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 7104 13268 7156 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 7288 13200 7340 13252
rect 9128 13200 9180 13252
rect 7196 13132 7248 13184
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 8668 13132 8720 13184
rect 9404 13200 9456 13252
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10416 13200 10468 13252
rect 10048 13132 10100 13184
rect 10600 13132 10652 13184
rect 12164 13132 12216 13184
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 13452 13268 13504 13320
rect 14464 13268 14516 13320
rect 16672 13268 16724 13320
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 14556 13200 14608 13252
rect 14740 13243 14792 13252
rect 14740 13209 14749 13243
rect 14749 13209 14783 13243
rect 14783 13209 14792 13243
rect 14740 13200 14792 13209
rect 16120 13200 16172 13252
rect 17408 13200 17460 13252
rect 13360 13132 13412 13184
rect 13636 13132 13688 13184
rect 15292 13132 15344 13184
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 16214 13030 16266 13082
rect 16278 13030 16330 13082
rect 16342 13030 16394 13082
rect 16406 13030 16458 13082
rect 16470 13030 16522 13082
rect 8668 12971 8720 12980
rect 8668 12937 8677 12971
rect 8677 12937 8711 12971
rect 8711 12937 8720 12971
rect 8668 12928 8720 12937
rect 9128 12928 9180 12980
rect 11060 12928 11112 12980
rect 4620 12860 4672 12912
rect 7748 12860 7800 12912
rect 9404 12860 9456 12912
rect 10140 12860 10192 12912
rect 12256 12928 12308 12980
rect 13176 12928 13228 12980
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 15476 12928 15528 12980
rect 16764 12928 16816 12980
rect 12164 12903 12216 12912
rect 12164 12869 12173 12903
rect 12173 12869 12207 12903
rect 12207 12869 12216 12903
rect 12164 12860 12216 12869
rect 14372 12860 14424 12912
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 3884 12835 3936 12844
rect 3884 12801 3893 12835
rect 3893 12801 3927 12835
rect 3927 12801 3936 12835
rect 3884 12792 3936 12801
rect 4068 12724 4120 12776
rect 6920 12792 6972 12844
rect 8116 12792 8168 12844
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 10232 12792 10284 12844
rect 10600 12792 10652 12844
rect 9220 12724 9272 12776
rect 10416 12724 10468 12776
rect 10968 12792 11020 12844
rect 14464 12792 14516 12844
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 15292 12792 15344 12844
rect 15936 12835 15988 12844
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 16672 12860 16724 12912
rect 17684 12860 17736 12912
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 18052 12835 18104 12844
rect 18052 12801 18070 12835
rect 18070 12801 18104 12835
rect 11152 12724 11204 12776
rect 12716 12724 12768 12776
rect 4804 12656 4856 12708
rect 7748 12656 7800 12708
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 14096 12724 14148 12776
rect 14556 12724 14608 12776
rect 16120 12724 16172 12776
rect 18052 12792 18104 12801
rect 15476 12588 15528 12640
rect 18236 12588 18288 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 3240 12384 3292 12436
rect 9864 12384 9916 12436
rect 2872 12316 2924 12368
rect 3148 12316 3200 12368
rect 3608 12316 3660 12368
rect 4620 12359 4672 12368
rect 4620 12325 4629 12359
rect 4629 12325 4663 12359
rect 4663 12325 4672 12359
rect 4620 12316 4672 12325
rect 7748 12359 7800 12368
rect 7748 12325 7757 12359
rect 7757 12325 7791 12359
rect 7791 12325 7800 12359
rect 7748 12316 7800 12325
rect 7932 12316 7984 12368
rect 13084 12384 13136 12436
rect 13176 12427 13228 12436
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 13360 12384 13412 12436
rect 14740 12384 14792 12436
rect 17408 12384 17460 12436
rect 17684 12427 17736 12436
rect 17684 12393 17693 12427
rect 17693 12393 17727 12427
rect 17727 12393 17736 12427
rect 17684 12384 17736 12393
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 2228 12112 2280 12164
rect 3884 12248 3936 12300
rect 6920 12248 6972 12300
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 3516 12180 3568 12189
rect 4804 12180 4856 12232
rect 3884 12112 3936 12164
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 7932 12112 7984 12164
rect 8852 12180 8904 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 10140 12180 10192 12232
rect 10324 12180 10376 12232
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 11152 12180 11204 12232
rect 11520 12180 11572 12232
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 18788 12316 18840 12368
rect 17592 12248 17644 12300
rect 14096 12180 14148 12232
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 14832 12180 14884 12232
rect 10416 12112 10468 12164
rect 10784 12112 10836 12164
rect 11796 12112 11848 12164
rect 14372 12112 14424 12164
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 16120 12180 16172 12232
rect 16764 12180 16816 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 17408 12180 17460 12232
rect 1492 12044 1544 12096
rect 2136 12044 2188 12096
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 6552 12044 6604 12096
rect 8024 12044 8076 12096
rect 8668 12044 8720 12096
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 9404 12044 9456 12096
rect 10324 12044 10376 12096
rect 11152 12044 11204 12096
rect 12716 12044 12768 12096
rect 14556 12087 14608 12096
rect 14556 12053 14565 12087
rect 14565 12053 14599 12087
rect 14599 12053 14608 12087
rect 14556 12044 14608 12053
rect 17408 12044 17460 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 16214 11942 16266 11994
rect 16278 11942 16330 11994
rect 16342 11942 16394 11994
rect 16406 11942 16458 11994
rect 16470 11942 16522 11994
rect 3424 11840 3476 11892
rect 6644 11840 6696 11892
rect 7196 11840 7248 11892
rect 8024 11883 8076 11892
rect 8024 11849 8033 11883
rect 8033 11849 8067 11883
rect 8067 11849 8076 11883
rect 8024 11840 8076 11849
rect 3700 11772 3752 11824
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 4620 11704 4672 11756
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 5816 11704 5868 11756
rect 7472 11704 7524 11756
rect 10048 11840 10100 11892
rect 10324 11840 10376 11892
rect 10968 11840 11020 11892
rect 8760 11772 8812 11824
rect 11888 11772 11940 11824
rect 13452 11772 13504 11824
rect 8576 11704 8628 11756
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 7932 11636 7984 11688
rect 8484 11636 8536 11688
rect 9036 11704 9088 11756
rect 8944 11679 8996 11688
rect 8944 11645 8953 11679
rect 8953 11645 8987 11679
rect 8987 11645 8996 11679
rect 8944 11636 8996 11645
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 10232 11747 10284 11756
rect 10232 11713 10241 11747
rect 10241 11713 10275 11747
rect 10275 11713 10284 11747
rect 10232 11704 10284 11713
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10600 11704 10652 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 10140 11636 10192 11688
rect 11520 11704 11572 11756
rect 12072 11704 12124 11756
rect 12532 11747 12584 11756
rect 12532 11713 12541 11747
rect 12541 11713 12575 11747
rect 12575 11713 12584 11747
rect 12532 11704 12584 11713
rect 12900 11704 12952 11756
rect 12992 11704 13044 11756
rect 14556 11840 14608 11892
rect 14832 11883 14884 11892
rect 14832 11849 14841 11883
rect 14841 11849 14875 11883
rect 14875 11849 14884 11883
rect 14832 11840 14884 11849
rect 14188 11704 14240 11756
rect 6552 11568 6604 11620
rect 11980 11636 12032 11688
rect 2228 11500 2280 11552
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 4068 11500 4120 11552
rect 8116 11500 8168 11552
rect 10600 11500 10652 11552
rect 10876 11500 10928 11552
rect 13820 11568 13872 11620
rect 14004 11679 14056 11688
rect 14004 11645 14013 11679
rect 14013 11645 14047 11679
rect 14047 11645 14056 11679
rect 15200 11704 15252 11756
rect 14004 11636 14056 11645
rect 17224 11704 17276 11756
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 13544 11500 13596 11552
rect 14372 11500 14424 11552
rect 15200 11500 15252 11552
rect 15568 11500 15620 11552
rect 15936 11500 15988 11552
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 18144 11500 18196 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 5080 11296 5132 11348
rect 6736 11296 6788 11348
rect 8760 11296 8812 11348
rect 4712 11228 4764 11280
rect 11704 11296 11756 11348
rect 12624 11296 12676 11348
rect 13176 11296 13228 11348
rect 13360 11296 13412 11348
rect 1492 11160 1544 11212
rect 7748 11160 7800 11212
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 9128 11160 9180 11212
rect 9312 11160 9364 11212
rect 9588 11160 9640 11212
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3516 11135 3568 11144
rect 3516 11101 3525 11135
rect 3525 11101 3559 11135
rect 3559 11101 3568 11135
rect 3516 11092 3568 11101
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 5816 11092 5868 11144
rect 6552 11092 6604 11144
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 8024 11092 8076 11144
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 2320 11067 2372 11076
rect 2320 11033 2329 11067
rect 2329 11033 2363 11067
rect 2363 11033 2372 11067
rect 2320 11024 2372 11033
rect 3424 11067 3476 11076
rect 3424 11033 3433 11067
rect 3433 11033 3467 11067
rect 3467 11033 3476 11067
rect 3424 11024 3476 11033
rect 7012 11024 7064 11076
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 9496 11024 9548 11076
rect 5540 10956 5592 11008
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 8944 10956 8996 11008
rect 10692 11160 10744 11212
rect 15476 11228 15528 11280
rect 16028 11228 16080 11280
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 9956 11135 10008 11144
rect 9956 11101 9965 11135
rect 9965 11101 9999 11135
rect 9999 11101 10008 11135
rect 9956 11092 10008 11101
rect 10416 11092 10468 11144
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 13084 11160 13136 11212
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 11796 11092 11848 11144
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 12440 11092 12492 11144
rect 14740 11135 14792 11144
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 15292 11160 15344 11212
rect 17316 11296 17368 11348
rect 16212 11228 16264 11280
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 16304 11092 16356 11144
rect 11612 11024 11664 11076
rect 11060 10956 11112 11008
rect 11336 10956 11388 11008
rect 11796 10956 11848 11008
rect 12900 10956 12952 11008
rect 13268 10999 13320 11008
rect 13636 11024 13688 11076
rect 13268 10965 13293 10999
rect 13293 10965 13320 10999
rect 13268 10956 13320 10965
rect 15844 11024 15896 11076
rect 16120 11024 16172 11076
rect 17408 11092 17460 11144
rect 18052 11024 18104 11076
rect 15200 10956 15252 11008
rect 15660 10956 15712 11008
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 16214 10854 16266 10906
rect 16278 10854 16330 10906
rect 16342 10854 16394 10906
rect 16406 10854 16458 10906
rect 16470 10854 16522 10906
rect 2320 10752 2372 10804
rect 3424 10752 3476 10804
rect 3884 10752 3936 10804
rect 5540 10684 5592 10736
rect 8116 10752 8168 10804
rect 9772 10752 9824 10804
rect 9956 10752 10008 10804
rect 10232 10752 10284 10804
rect 10508 10752 10560 10804
rect 10600 10752 10652 10804
rect 11980 10752 12032 10804
rect 12808 10795 12860 10804
rect 12808 10761 12817 10795
rect 12817 10761 12851 10795
rect 12851 10761 12860 10795
rect 12808 10752 12860 10761
rect 14740 10752 14792 10804
rect 3332 10616 3384 10668
rect 4160 10616 4212 10668
rect 5080 10616 5132 10668
rect 5908 10616 5960 10668
rect 2964 10548 3016 10600
rect 4804 10548 4856 10600
rect 6644 10616 6696 10668
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7656 10659 7708 10668
rect 7656 10625 7667 10659
rect 7667 10625 7708 10659
rect 7656 10616 7708 10625
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 8116 10616 8168 10668
rect 9864 10684 9916 10736
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9496 10616 9548 10668
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 10508 10616 10560 10668
rect 11336 10684 11388 10736
rect 7472 10548 7524 10600
rect 8852 10548 8904 10600
rect 11612 10616 11664 10668
rect 3976 10480 4028 10532
rect 10140 10480 10192 10532
rect 10416 10480 10468 10532
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 14832 10684 14884 10736
rect 15660 10752 15712 10804
rect 17960 10752 18012 10804
rect 15200 10727 15252 10736
rect 15200 10693 15210 10727
rect 15210 10693 15244 10727
rect 15244 10693 15252 10727
rect 15200 10684 15252 10693
rect 15384 10684 15436 10736
rect 15476 10684 15528 10736
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 11888 10548 11940 10600
rect 12808 10616 12860 10668
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 13912 10616 13964 10668
rect 14280 10616 14332 10668
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 18144 10727 18196 10736
rect 18144 10693 18153 10727
rect 18153 10693 18187 10727
rect 18187 10693 18196 10727
rect 18144 10684 18196 10693
rect 18236 10727 18288 10736
rect 18236 10693 18245 10727
rect 18245 10693 18279 10727
rect 18279 10693 18288 10727
rect 18236 10684 18288 10693
rect 12532 10548 12584 10600
rect 13636 10548 13688 10600
rect 14924 10548 14976 10600
rect 17224 10616 17276 10668
rect 15200 10548 15252 10600
rect 15936 10548 15988 10600
rect 16764 10548 16816 10600
rect 4712 10412 4764 10464
rect 5540 10412 5592 10464
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 8392 10412 8444 10464
rect 12624 10480 12676 10532
rect 13084 10480 13136 10532
rect 13268 10480 13320 10532
rect 11152 10412 11204 10464
rect 12256 10412 12308 10464
rect 12716 10412 12768 10464
rect 13728 10412 13780 10464
rect 16120 10480 16172 10532
rect 17224 10523 17276 10532
rect 17224 10489 17233 10523
rect 17233 10489 17267 10523
rect 17267 10489 17276 10523
rect 17224 10480 17276 10489
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 7656 10140 7708 10192
rect 7932 10183 7984 10192
rect 7932 10149 7941 10183
rect 7941 10149 7975 10183
rect 7975 10149 7984 10183
rect 7932 10140 7984 10149
rect 2228 10004 2280 10056
rect 5540 10004 5592 10056
rect 5816 10004 5868 10056
rect 7380 10072 7432 10124
rect 8944 10208 8996 10260
rect 9312 10208 9364 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 10232 10208 10284 10260
rect 9772 10140 9824 10192
rect 10416 10140 10468 10192
rect 9036 10072 9088 10124
rect 8024 10004 8076 10056
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 8668 10004 8720 10056
rect 9220 10047 9272 10056
rect 9220 10013 9230 10047
rect 9230 10013 9264 10047
rect 9264 10013 9272 10047
rect 9220 10004 9272 10013
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 4620 9936 4672 9988
rect 4804 9936 4856 9988
rect 2044 9868 2096 9920
rect 5908 9868 5960 9920
rect 6184 9911 6236 9920
rect 6184 9877 6193 9911
rect 6193 9877 6227 9911
rect 6227 9877 6236 9911
rect 6184 9868 6236 9877
rect 7196 9868 7248 9920
rect 7564 9936 7616 9988
rect 8760 9868 8812 9920
rect 9404 9868 9456 9920
rect 9772 9936 9824 9988
rect 11888 10208 11940 10260
rect 12624 10208 12676 10260
rect 12716 10208 12768 10260
rect 15292 10251 15344 10260
rect 15292 10217 15301 10251
rect 15301 10217 15335 10251
rect 15335 10217 15344 10251
rect 15292 10208 15344 10217
rect 11428 10140 11480 10192
rect 10692 10004 10744 10056
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 12624 10072 12676 10124
rect 13084 10183 13136 10192
rect 13084 10149 13093 10183
rect 13093 10149 13127 10183
rect 13127 10149 13136 10183
rect 13084 10140 13136 10149
rect 11796 10004 11848 10056
rect 12900 10004 12952 10056
rect 13176 10004 13228 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 15016 10140 15068 10192
rect 17960 10140 18012 10192
rect 17040 10072 17092 10124
rect 10416 9936 10468 9988
rect 10508 9936 10560 9988
rect 9588 9868 9640 9920
rect 10600 9868 10652 9920
rect 12808 9936 12860 9988
rect 13820 10004 13872 10056
rect 15660 10004 15712 10056
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 18144 10004 18196 10056
rect 10876 9868 10928 9920
rect 11520 9911 11572 9920
rect 11520 9877 11529 9911
rect 11529 9877 11563 9911
rect 11563 9877 11572 9911
rect 11520 9868 11572 9877
rect 11612 9868 11664 9920
rect 14096 9936 14148 9988
rect 14832 9936 14884 9988
rect 13084 9868 13136 9920
rect 13912 9868 13964 9920
rect 17408 9936 17460 9988
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 16214 9766 16266 9818
rect 16278 9766 16330 9818
rect 16342 9766 16394 9818
rect 16406 9766 16458 9818
rect 16470 9766 16522 9818
rect 5908 9707 5960 9716
rect 5908 9673 5917 9707
rect 5917 9673 5951 9707
rect 5951 9673 5960 9707
rect 5908 9664 5960 9673
rect 7472 9707 7524 9716
rect 7472 9673 7481 9707
rect 7481 9673 7515 9707
rect 7515 9673 7524 9707
rect 7472 9664 7524 9673
rect 7564 9664 7616 9716
rect 8668 9664 8720 9716
rect 9404 9664 9456 9716
rect 9956 9664 10008 9716
rect 12072 9664 12124 9716
rect 9220 9596 9272 9648
rect 10692 9639 10744 9648
rect 2228 9528 2280 9580
rect 3056 9528 3108 9580
rect 4988 9528 5040 9580
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 7932 9528 7984 9580
rect 9036 9571 9088 9580
rect 9036 9537 9045 9571
rect 9045 9537 9079 9571
rect 9079 9537 9088 9571
rect 9036 9528 9088 9537
rect 10692 9605 10701 9639
rect 10701 9605 10735 9639
rect 10735 9605 10744 9639
rect 10692 9596 10744 9605
rect 1860 9392 1912 9444
rect 4620 9392 4672 9444
rect 5816 9460 5868 9512
rect 7656 9460 7708 9512
rect 8576 9460 8628 9512
rect 9404 9571 9456 9580
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 9404 9528 9456 9537
rect 9588 9528 9640 9580
rect 12900 9664 12952 9716
rect 13728 9664 13780 9716
rect 14556 9664 14608 9716
rect 15292 9664 15344 9716
rect 11704 9528 11756 9580
rect 12716 9596 12768 9648
rect 13084 9596 13136 9648
rect 14096 9596 14148 9648
rect 14188 9639 14240 9648
rect 14188 9605 14197 9639
rect 14197 9605 14231 9639
rect 14231 9605 14240 9639
rect 14188 9596 14240 9605
rect 14464 9596 14516 9648
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 12072 9460 12124 9512
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 12992 9528 13044 9580
rect 13360 9528 13412 9580
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 15476 9596 15528 9648
rect 16764 9596 16816 9648
rect 15108 9528 15160 9580
rect 15200 9528 15252 9580
rect 17132 9528 17184 9580
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 6552 9392 6604 9444
rect 7564 9392 7616 9444
rect 3240 9324 3292 9376
rect 6828 9324 6880 9376
rect 8944 9324 8996 9376
rect 10140 9392 10192 9444
rect 11888 9392 11940 9444
rect 13360 9392 13412 9444
rect 13452 9392 13504 9444
rect 13636 9392 13688 9444
rect 14924 9392 14976 9444
rect 11612 9324 11664 9376
rect 15752 9392 15804 9444
rect 15936 9392 15988 9444
rect 17592 9324 17644 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 3056 9163 3108 9172
rect 3056 9129 3065 9163
rect 3065 9129 3099 9163
rect 3099 9129 3108 9163
rect 3056 9120 3108 9129
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 7196 9120 7248 9172
rect 9404 9120 9456 9172
rect 9864 9120 9916 9172
rect 1308 8984 1360 9036
rect 4620 9052 4672 9104
rect 1216 8916 1268 8968
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 2136 8916 2188 8968
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4712 8984 4764 9036
rect 6092 8916 6144 8968
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 9680 9052 9732 9104
rect 7288 9027 7340 9036
rect 7288 8993 7297 9027
rect 7297 8993 7331 9027
rect 7331 8993 7340 9027
rect 7288 8984 7340 8993
rect 7932 8984 7984 9036
rect 4896 8891 4948 8900
rect 4896 8857 4905 8891
rect 4905 8857 4939 8891
rect 4939 8857 4948 8891
rect 4896 8848 4948 8857
rect 6368 8891 6420 8900
rect 6368 8857 6377 8891
rect 6377 8857 6411 8891
rect 6411 8857 6420 8891
rect 6368 8848 6420 8857
rect 6920 8891 6972 8900
rect 6920 8857 6929 8891
rect 6929 8857 6963 8891
rect 6963 8857 6972 8891
rect 6920 8848 6972 8857
rect 2964 8780 3016 8832
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 5540 8780 5592 8832
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 7104 8780 7156 8832
rect 7380 8959 7432 8968
rect 9496 8984 9548 9036
rect 11704 9120 11756 9172
rect 12992 9120 13044 9172
rect 13636 9052 13688 9104
rect 7380 8925 7401 8959
rect 7401 8925 7432 8959
rect 7380 8916 7432 8925
rect 7840 8891 7892 8900
rect 7840 8857 7849 8891
rect 7849 8857 7883 8891
rect 7883 8857 7892 8891
rect 7840 8848 7892 8857
rect 8760 8848 8812 8900
rect 7656 8780 7708 8832
rect 9772 8916 9824 8968
rect 9956 8916 10008 8968
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 10876 8984 10928 9036
rect 12532 9027 12584 9036
rect 10232 8848 10284 8900
rect 10692 8916 10744 8968
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 14464 9052 14516 9104
rect 14832 9052 14884 9104
rect 10784 8891 10836 8900
rect 10784 8857 10793 8891
rect 10793 8857 10827 8891
rect 10827 8857 10836 8891
rect 10784 8848 10836 8857
rect 11704 8916 11756 8968
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 12900 8959 12952 8968
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 13268 8916 13320 8968
rect 13452 8916 13504 8968
rect 14556 8984 14608 9036
rect 11980 8891 12032 8900
rect 11980 8857 11989 8891
rect 11989 8857 12023 8891
rect 12023 8857 12032 8891
rect 11980 8848 12032 8857
rect 10692 8780 10744 8832
rect 10968 8780 11020 8832
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 15384 9120 15436 9172
rect 17224 9120 17276 9172
rect 15384 8916 15436 8968
rect 15476 8916 15528 8968
rect 17592 9095 17644 9104
rect 17592 9061 17601 9095
rect 17601 9061 17635 9095
rect 17635 9061 17644 9095
rect 17592 9052 17644 9061
rect 16764 8916 16816 8968
rect 17408 8984 17460 9036
rect 17132 8959 17184 8968
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 17960 8959 18012 8968
rect 17960 8925 18004 8959
rect 18004 8925 18012 8959
rect 17960 8916 18012 8925
rect 15752 8848 15804 8900
rect 13084 8780 13136 8832
rect 13360 8780 13412 8832
rect 14280 8780 14332 8832
rect 15844 8780 15896 8832
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 16214 8678 16266 8730
rect 16278 8678 16330 8730
rect 16342 8678 16394 8730
rect 16406 8678 16458 8730
rect 16470 8678 16522 8730
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 7288 8576 7340 8628
rect 7564 8576 7616 8628
rect 13268 8576 13320 8628
rect 14372 8576 14424 8628
rect 14556 8576 14608 8628
rect 15200 8576 15252 8628
rect 15844 8619 15896 8628
rect 15844 8585 15853 8619
rect 15853 8585 15887 8619
rect 15887 8585 15896 8619
rect 15844 8576 15896 8585
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 6460 8508 6512 8560
rect 6184 8440 6236 8492
rect 7012 8508 7064 8560
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 8024 8508 8076 8560
rect 9772 8551 9824 8560
rect 9772 8517 9781 8551
rect 9781 8517 9815 8551
rect 9815 8517 9824 8551
rect 9772 8508 9824 8517
rect 10232 8508 10284 8560
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 3516 8372 3568 8424
rect 6368 8372 6420 8424
rect 4896 8304 4948 8356
rect 7104 8347 7156 8356
rect 7104 8313 7113 8347
rect 7113 8313 7147 8347
rect 7147 8313 7156 8347
rect 7104 8304 7156 8313
rect 7472 8372 7524 8424
rect 8116 8440 8168 8492
rect 8576 8440 8628 8492
rect 9312 8440 9364 8492
rect 9588 8483 9640 8492
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 12072 8508 12124 8560
rect 13544 8508 13596 8560
rect 10048 8440 10100 8449
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 11060 8440 11112 8492
rect 11428 8440 11480 8492
rect 9864 8372 9916 8424
rect 11888 8372 11940 8424
rect 12716 8440 12768 8492
rect 9496 8304 9548 8356
rect 2228 8236 2280 8288
rect 8392 8236 8444 8288
rect 8576 8236 8628 8288
rect 9772 8254 9824 8306
rect 10140 8304 10192 8356
rect 10692 8304 10744 8356
rect 10968 8304 11020 8356
rect 12072 8304 12124 8356
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13360 8440 13412 8492
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 14464 8440 14516 8492
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 10416 8236 10468 8288
rect 11796 8236 11848 8288
rect 13452 8304 13504 8356
rect 13820 8304 13872 8356
rect 13268 8236 13320 8288
rect 13912 8236 13964 8288
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 16948 8576 17000 8628
rect 17592 8508 17644 8560
rect 16672 8372 16724 8424
rect 17776 8304 17828 8356
rect 14648 8279 14700 8288
rect 14648 8245 14657 8279
rect 14657 8245 14691 8279
rect 14691 8245 14700 8279
rect 14648 8236 14700 8245
rect 15936 8236 15988 8288
rect 16580 8236 16632 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 3608 8032 3660 8084
rect 6092 8032 6144 8084
rect 9496 8032 9548 8084
rect 11244 8032 11296 8084
rect 2964 7896 3016 7948
rect 4896 7964 4948 8016
rect 6920 7964 6972 8016
rect 9312 7964 9364 8016
rect 12716 8032 12768 8084
rect 5540 7896 5592 7948
rect 6184 7896 6236 7948
rect 6460 7896 6512 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 2596 7828 2648 7880
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 7104 7896 7156 7948
rect 8024 7896 8076 7948
rect 8300 7896 8352 7948
rect 9956 7896 10008 7948
rect 10416 7896 10468 7948
rect 12072 7896 12124 7948
rect 12900 7964 12952 8016
rect 3884 7760 3936 7812
rect 7564 7828 7616 7880
rect 7748 7828 7800 7880
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 8392 7828 8444 7880
rect 10140 7828 10192 7880
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 10508 7760 10560 7812
rect 11796 7828 11848 7880
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 15476 7964 15528 8016
rect 15752 7964 15804 8016
rect 13912 7896 13964 7948
rect 14740 7939 14792 7948
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 16028 7896 16080 7948
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 14372 7871 14424 7880
rect 14372 7837 14381 7871
rect 14381 7837 14415 7871
rect 14415 7837 14424 7871
rect 14372 7828 14424 7837
rect 14648 7828 14700 7880
rect 15016 7828 15068 7880
rect 16580 7828 16632 7880
rect 16856 7871 16908 7880
rect 16856 7837 16865 7871
rect 16865 7837 16899 7871
rect 16899 7837 16908 7871
rect 16856 7828 16908 7837
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 18328 7828 18380 7880
rect 12808 7760 12860 7812
rect 13176 7760 13228 7812
rect 16212 7803 16264 7812
rect 16212 7769 16221 7803
rect 16221 7769 16255 7803
rect 16255 7769 16264 7803
rect 16212 7760 16264 7769
rect 16948 7760 17000 7812
rect 6736 7692 6788 7744
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 7840 7692 7892 7744
rect 9680 7692 9732 7744
rect 12716 7692 12768 7744
rect 18144 7692 18196 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 16214 7590 16266 7642
rect 16278 7590 16330 7642
rect 16342 7590 16394 7642
rect 16406 7590 16458 7642
rect 16470 7590 16522 7642
rect 2688 7488 2740 7540
rect 8116 7488 8168 7540
rect 10232 7488 10284 7540
rect 10968 7488 11020 7540
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2136 7352 2188 7404
rect 2412 7395 2464 7404
rect 2412 7361 2421 7395
rect 2421 7361 2455 7395
rect 2455 7361 2464 7395
rect 2412 7352 2464 7361
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 2688 7352 2740 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 6368 7420 6420 7472
rect 6736 7420 6788 7472
rect 2320 7216 2372 7268
rect 2596 7148 2648 7200
rect 2780 7216 2832 7268
rect 4804 7284 4856 7336
rect 7104 7216 7156 7268
rect 9588 7420 9640 7472
rect 10416 7420 10468 7472
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 16764 7531 16816 7540
rect 16764 7497 16773 7531
rect 16773 7497 16807 7531
rect 16807 7497 16816 7531
rect 16764 7488 16816 7497
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 8116 7352 8168 7404
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 9312 7352 9364 7404
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 13728 7420 13780 7472
rect 10048 7284 10100 7336
rect 8760 7216 8812 7268
rect 11888 7216 11940 7268
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 8484 7148 8536 7200
rect 13452 7352 13504 7404
rect 15476 7420 15528 7472
rect 15936 7463 15988 7472
rect 15936 7429 15945 7463
rect 15945 7429 15979 7463
rect 15979 7429 15988 7463
rect 15936 7420 15988 7429
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 16028 7352 16080 7404
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 12992 7327 13044 7336
rect 12992 7293 13001 7327
rect 13001 7293 13035 7327
rect 13035 7293 13044 7327
rect 12992 7284 13044 7293
rect 13268 7284 13320 7336
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 16856 7284 16908 7336
rect 14280 7259 14332 7268
rect 14280 7225 14289 7259
rect 14289 7225 14323 7259
rect 14323 7225 14332 7259
rect 14280 7216 14332 7225
rect 15108 7259 15160 7268
rect 15108 7225 15117 7259
rect 15117 7225 15151 7259
rect 15151 7225 15160 7259
rect 15108 7216 15160 7225
rect 15752 7148 15804 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 2412 6944 2464 6996
rect 2780 6944 2832 6996
rect 1676 6876 1728 6928
rect 3424 6944 3476 6996
rect 4068 6944 4120 6996
rect 4988 6944 5040 6996
rect 17040 6944 17092 6996
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 2320 6740 2372 6792
rect 2504 6783 2556 6792
rect 2504 6749 2513 6783
rect 2513 6749 2547 6783
rect 2547 6749 2556 6783
rect 2504 6740 2556 6749
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 2872 6672 2924 6724
rect 2136 6604 2188 6656
rect 3608 6604 3660 6656
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 6736 6851 6788 6860
rect 6736 6817 6745 6851
rect 6745 6817 6779 6851
rect 6779 6817 6788 6851
rect 6736 6808 6788 6817
rect 6828 6740 6880 6792
rect 7012 6876 7064 6928
rect 8116 6919 8168 6928
rect 8116 6885 8125 6919
rect 8125 6885 8159 6919
rect 8159 6885 8168 6919
rect 8116 6876 8168 6885
rect 9588 6808 9640 6860
rect 10876 6876 10928 6928
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 8760 6672 8812 6724
rect 11060 6740 11112 6792
rect 13084 6876 13136 6928
rect 14280 6808 14332 6860
rect 14832 6851 14884 6860
rect 14832 6817 14841 6851
rect 14841 6817 14875 6851
rect 14875 6817 14884 6851
rect 14832 6808 14884 6817
rect 12716 6783 12768 6792
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 10048 6672 10100 6724
rect 8024 6604 8076 6656
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 9680 6604 9732 6656
rect 12072 6672 12124 6724
rect 12900 6740 12952 6792
rect 13360 6740 13412 6792
rect 15200 6783 15252 6792
rect 15200 6749 15209 6783
rect 15209 6749 15243 6783
rect 15243 6749 15252 6783
rect 15200 6740 15252 6749
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 16120 6740 16172 6792
rect 16580 6740 16632 6792
rect 16856 6740 16908 6792
rect 11060 6604 11112 6656
rect 15476 6672 15528 6724
rect 12808 6604 12860 6656
rect 14464 6604 14516 6656
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 14648 6604 14700 6656
rect 15568 6604 15620 6656
rect 15752 6604 15804 6656
rect 17316 6740 17368 6792
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 18328 6604 18380 6656
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 16214 6502 16266 6554
rect 16278 6502 16330 6554
rect 16342 6502 16394 6554
rect 16406 6502 16458 6554
rect 16470 6502 16522 6554
rect 2228 6400 2280 6452
rect 2504 6400 2556 6452
rect 3240 6400 3292 6452
rect 2412 6332 2464 6384
rect 1768 6264 1820 6316
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 3240 6307 3292 6316
rect 1860 6196 1912 6248
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 2228 6128 2280 6180
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 6736 6400 6788 6452
rect 10508 6400 10560 6452
rect 10784 6400 10836 6452
rect 14740 6400 14792 6452
rect 17316 6400 17368 6452
rect 4896 6264 4948 6316
rect 6644 6264 6696 6316
rect 8576 6264 8628 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 10048 6332 10100 6384
rect 3332 6060 3384 6112
rect 3976 6060 4028 6112
rect 6736 6128 6788 6180
rect 8116 6196 8168 6248
rect 9864 6264 9916 6316
rect 10140 6264 10192 6316
rect 13268 6332 13320 6384
rect 14648 6332 14700 6384
rect 15108 6332 15160 6384
rect 17776 6332 17828 6384
rect 11244 6264 11296 6316
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16028 6307 16080 6316
rect 16028 6273 16037 6307
rect 16037 6273 16071 6307
rect 16071 6273 16080 6307
rect 16028 6264 16080 6273
rect 8760 6128 8812 6180
rect 9588 6128 9640 6180
rect 13360 6196 13412 6248
rect 14832 6196 14884 6248
rect 17316 6307 17368 6316
rect 17316 6273 17325 6307
rect 17325 6273 17359 6307
rect 17359 6273 17368 6307
rect 17316 6264 17368 6273
rect 10324 6128 10376 6180
rect 4620 6060 4672 6112
rect 5448 6060 5500 6112
rect 6092 6060 6144 6112
rect 7104 6060 7156 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 14004 6128 14056 6180
rect 15936 6128 15988 6180
rect 18328 6128 18380 6180
rect 12992 6060 13044 6112
rect 13912 6103 13964 6112
rect 13912 6069 13921 6103
rect 13921 6069 13955 6103
rect 13955 6069 13964 6103
rect 13912 6060 13964 6069
rect 14372 6060 14424 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 4436 5856 4488 5908
rect 4804 5856 4856 5908
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 9588 5856 9640 5908
rect 12716 5856 12768 5908
rect 13360 5856 13412 5908
rect 16028 5856 16080 5908
rect 18420 5856 18472 5908
rect 3332 5788 3384 5840
rect 3148 5720 3200 5772
rect 5356 5788 5408 5840
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 2964 5652 3016 5704
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3332 5584 3384 5636
rect 6092 5720 6144 5772
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 4436 5652 4488 5704
rect 4988 5695 5040 5704
rect 4988 5661 4997 5695
rect 4997 5661 5031 5695
rect 5031 5661 5040 5695
rect 4988 5652 5040 5661
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 6000 5652 6052 5704
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 9128 5652 9180 5704
rect 5080 5584 5132 5636
rect 8116 5584 8168 5636
rect 9864 5652 9916 5704
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 11980 5720 12032 5772
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 12624 5695 12676 5704
rect 12624 5661 12633 5695
rect 12633 5661 12667 5695
rect 12667 5661 12676 5695
rect 12624 5652 12676 5661
rect 12900 5652 12952 5704
rect 13084 5652 13136 5704
rect 13360 5695 13412 5704
rect 13360 5661 13369 5695
rect 13369 5661 13403 5695
rect 13403 5661 13412 5695
rect 13360 5652 13412 5661
rect 13912 5720 13964 5772
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 14556 5720 14608 5772
rect 16120 5720 16172 5772
rect 16580 5720 16632 5772
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 17776 5652 17828 5704
rect 11612 5584 11664 5636
rect 14096 5584 14148 5636
rect 16856 5584 16908 5636
rect 4712 5516 4764 5568
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 9680 5516 9732 5568
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 16214 5414 16266 5466
rect 16278 5414 16330 5466
rect 16342 5414 16394 5466
rect 16406 5414 16458 5466
rect 16470 5414 16522 5466
rect 2228 5312 2280 5364
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 940 5176 992 5228
rect 4712 5287 4764 5296
rect 4712 5253 4721 5287
rect 4721 5253 4755 5287
rect 4755 5253 4764 5287
rect 4712 5244 4764 5253
rect 4804 5244 4856 5296
rect 4988 5312 5040 5364
rect 6000 5355 6052 5364
rect 6000 5321 6009 5355
rect 6009 5321 6043 5355
rect 6043 5321 6052 5355
rect 6000 5312 6052 5321
rect 8116 5312 8168 5364
rect 8852 5312 8904 5364
rect 3056 5176 3108 5228
rect 3148 5219 3200 5228
rect 3148 5185 3157 5219
rect 3157 5185 3191 5219
rect 3191 5185 3200 5219
rect 3148 5176 3200 5185
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 4620 5176 4672 5228
rect 2964 5108 3016 5160
rect 5080 5176 5132 5228
rect 5448 5176 5500 5228
rect 5356 5108 5408 5160
rect 6736 5176 6788 5228
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 6644 5108 6696 5160
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 7104 5108 7156 5160
rect 9128 5244 9180 5296
rect 5172 5040 5224 5092
rect 6552 5040 6604 5092
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 8208 5108 8260 5160
rect 8760 5176 8812 5228
rect 9864 5312 9916 5364
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 13176 5312 13228 5364
rect 15476 5355 15528 5364
rect 15476 5321 15485 5355
rect 15485 5321 15519 5355
rect 15519 5321 15528 5355
rect 15476 5312 15528 5321
rect 16120 5312 16172 5364
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 17224 5355 17276 5364
rect 17224 5321 17233 5355
rect 17233 5321 17267 5355
rect 17267 5321 17276 5355
rect 17224 5312 17276 5321
rect 9312 5244 9364 5296
rect 9680 5244 9732 5296
rect 11888 5287 11940 5296
rect 11888 5253 11897 5287
rect 11897 5253 11931 5287
rect 11931 5253 11940 5287
rect 11888 5244 11940 5253
rect 12624 5244 12676 5296
rect 11612 5219 11664 5228
rect 11612 5185 11621 5219
rect 11621 5185 11655 5219
rect 11655 5185 11664 5219
rect 11612 5176 11664 5185
rect 13912 5244 13964 5296
rect 14004 5287 14056 5296
rect 14004 5253 14013 5287
rect 14013 5253 14047 5287
rect 14047 5253 14056 5287
rect 14004 5244 14056 5253
rect 14096 5244 14148 5296
rect 15844 5176 15896 5228
rect 16120 5176 16172 5228
rect 16672 5176 16724 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 8944 5108 8996 5160
rect 13084 5108 13136 5160
rect 9772 4972 9824 5024
rect 16028 5015 16080 5024
rect 16028 4981 16037 5015
rect 16037 4981 16071 5015
rect 16071 4981 16080 5015
rect 16028 4972 16080 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 6644 4768 6696 4820
rect 7564 4768 7616 4820
rect 8944 4768 8996 4820
rect 9864 4768 9916 4820
rect 11152 4768 11204 4820
rect 11612 4768 11664 4820
rect 12624 4768 12676 4820
rect 4804 4700 4856 4752
rect 7012 4700 7064 4752
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 1952 4564 2004 4616
rect 3424 4564 3476 4616
rect 6460 4632 6512 4684
rect 6644 4632 6696 4684
rect 6920 4632 6972 4684
rect 5172 4564 5224 4616
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 8668 4632 8720 4684
rect 8208 4564 8260 4616
rect 8944 4564 8996 4616
rect 12440 4632 12492 4684
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 3608 4496 3660 4548
rect 1860 4428 1912 4480
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 4528 4496 4580 4548
rect 5264 4496 5316 4548
rect 4712 4428 4764 4480
rect 6920 4428 6972 4480
rect 7564 4471 7616 4480
rect 7564 4437 7573 4471
rect 7573 4437 7607 4471
rect 7607 4437 7616 4471
rect 7564 4428 7616 4437
rect 9772 4496 9824 4548
rect 13084 4768 13136 4820
rect 13912 4811 13964 4820
rect 13912 4777 13921 4811
rect 13921 4777 13955 4811
rect 13955 4777 13964 4811
rect 13912 4768 13964 4777
rect 15200 4768 15252 4820
rect 14372 4496 14424 4548
rect 16028 4496 16080 4548
rect 12440 4428 12492 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 16214 4326 16266 4378
rect 16278 4326 16330 4378
rect 16342 4326 16394 4378
rect 16406 4326 16458 4378
rect 16470 4326 16522 4378
rect 3424 4224 3476 4276
rect 2780 4199 2832 4208
rect 2780 4165 2789 4199
rect 2789 4165 2823 4199
rect 2823 4165 2832 4199
rect 2780 4156 2832 4165
rect 1768 4088 1820 4140
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 2320 4088 2372 4140
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 4712 4131 4764 4140
rect 4712 4097 4721 4131
rect 4721 4097 4755 4131
rect 4755 4097 4764 4131
rect 4712 4088 4764 4097
rect 5632 4156 5684 4208
rect 6828 4156 6880 4208
rect 5172 3952 5224 4004
rect 6368 4020 6420 4072
rect 7012 4088 7064 4140
rect 7564 4156 7616 4208
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 9588 4088 9640 4140
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 7104 4020 7156 4072
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 8116 4020 8168 4072
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9404 4020 9456 4072
rect 9772 4020 9824 4072
rect 11888 4088 11940 4140
rect 13912 4224 13964 4276
rect 12440 4020 12492 4072
rect 13084 4020 13136 4072
rect 11152 3952 11204 4004
rect 12072 3952 12124 4004
rect 15844 4088 15896 4140
rect 16580 4088 16632 4140
rect 16948 4088 17000 4140
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 2964 3884 3016 3936
rect 8024 3884 8076 3936
rect 9772 3884 9824 3936
rect 9956 3884 10008 3936
rect 10784 3927 10836 3936
rect 10784 3893 10793 3927
rect 10793 3893 10827 3927
rect 10827 3893 10836 3927
rect 10784 3884 10836 3893
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 16672 3884 16724 3936
rect 17408 4063 17460 4072
rect 17408 4029 17417 4063
rect 17417 4029 17451 4063
rect 17451 4029 17460 4063
rect 17408 4020 17460 4029
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 2872 3680 2924 3732
rect 5080 3680 5132 3732
rect 7472 3680 7524 3732
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 1952 3612 2004 3664
rect 5356 3612 5408 3664
rect 10140 3680 10192 3732
rect 12072 3680 12124 3732
rect 1860 3544 1912 3596
rect 2320 3544 2372 3596
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 1308 3476 1360 3528
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 2044 3476 2096 3528
rect 4804 3476 4856 3528
rect 3700 3408 3752 3460
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 7748 3476 7800 3528
rect 9496 3612 9548 3664
rect 9956 3612 10008 3664
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 9404 3544 9456 3596
rect 14924 3680 14976 3732
rect 16580 3680 16632 3732
rect 17040 3723 17092 3732
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 1860 3340 1912 3392
rect 6736 3340 6788 3392
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 9956 3476 10008 3528
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 13912 3544 13964 3596
rect 17408 3544 17460 3596
rect 11796 3408 11848 3460
rect 12992 3340 13044 3392
rect 16028 3476 16080 3528
rect 16672 3476 16724 3528
rect 17132 3476 17184 3528
rect 16672 3383 16724 3392
rect 16672 3349 16681 3383
rect 16681 3349 16715 3383
rect 16715 3349 16724 3383
rect 16672 3340 16724 3349
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 16214 3238 16266 3290
rect 16278 3238 16330 3290
rect 16342 3238 16394 3290
rect 16406 3238 16458 3290
rect 16470 3238 16522 3290
rect 2320 3136 2372 3188
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 4712 3136 4764 3188
rect 2136 3000 2188 3052
rect 4804 3068 4856 3120
rect 5908 3136 5960 3188
rect 7748 3136 7800 3188
rect 9036 3136 9088 3188
rect 9588 3136 9640 3188
rect 9680 3136 9732 3188
rect 1308 2932 1360 2984
rect 2780 3000 2832 3052
rect 3424 3043 3476 3052
rect 3424 3009 3433 3043
rect 3433 3009 3467 3043
rect 3467 3009 3476 3043
rect 3424 3000 3476 3009
rect 4620 3000 4672 3052
rect 5448 3000 5500 3052
rect 6736 3068 6788 3120
rect 7840 3068 7892 3120
rect 8484 3111 8536 3120
rect 8484 3077 8493 3111
rect 8493 3077 8527 3111
rect 8527 3077 8536 3111
rect 8484 3068 8536 3077
rect 8668 3111 8720 3120
rect 8668 3077 8693 3111
rect 8693 3077 8720 3111
rect 13912 3136 13964 3188
rect 16672 3136 16724 3188
rect 8668 3068 8720 3077
rect 5080 2932 5132 2984
rect 12072 3068 12124 3120
rect 12992 3068 13044 3120
rect 9220 3000 9272 3052
rect 9772 3000 9824 3052
rect 11244 3000 11296 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 15568 3000 15620 3052
rect 15844 3000 15896 3052
rect 16580 3000 16632 3052
rect 17408 3000 17460 3052
rect 17684 3043 17736 3052
rect 17684 3009 17693 3043
rect 17693 3009 17727 3043
rect 17727 3009 17736 3043
rect 17684 3000 17736 3009
rect 8484 2864 8536 2916
rect 10232 2932 10284 2984
rect 10968 2864 11020 2916
rect 2136 2796 2188 2848
rect 3976 2796 4028 2848
rect 5264 2796 5316 2848
rect 7012 2796 7064 2848
rect 7196 2796 7248 2848
rect 7472 2839 7524 2848
rect 7472 2805 7481 2839
rect 7481 2805 7515 2839
rect 7515 2805 7524 2839
rect 7472 2796 7524 2805
rect 8300 2796 8352 2848
rect 8760 2796 8812 2848
rect 11152 2932 11204 2984
rect 12072 2932 12124 2984
rect 12072 2796 12124 2848
rect 16028 2796 16080 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 2044 2592 2096 2644
rect 2136 2592 2188 2644
rect 2780 2592 2832 2644
rect 5172 2592 5224 2644
rect 3424 2567 3476 2576
rect 3424 2533 3433 2567
rect 3433 2533 3467 2567
rect 3467 2533 3476 2567
rect 3424 2524 3476 2533
rect 1952 2456 2004 2508
rect 6000 2592 6052 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 6920 2592 6972 2644
rect 1860 2431 1912 2440
rect 1860 2397 1870 2431
rect 1870 2397 1904 2431
rect 1904 2397 1912 2431
rect 1860 2388 1912 2397
rect 2964 2388 3016 2440
rect 3700 2388 3752 2440
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 4712 2388 4764 2440
rect 5080 2388 5132 2440
rect 5540 2388 5592 2440
rect 5908 2388 5960 2440
rect 7472 2456 7524 2508
rect 8024 2456 8076 2508
rect 9864 2592 9916 2644
rect 10784 2592 10836 2644
rect 11244 2592 11296 2644
rect 12992 2635 13044 2644
rect 12992 2601 13001 2635
rect 13001 2601 13035 2635
rect 13035 2601 13044 2635
rect 12992 2592 13044 2601
rect 7012 2388 7064 2440
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 7564 2388 7616 2440
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 9680 2388 9732 2440
rect 10140 2456 10192 2508
rect 10232 2456 10284 2508
rect 17684 2524 17736 2576
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 15568 2456 15620 2508
rect 15752 2499 15804 2508
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 15752 2456 15804 2465
rect 7840 2363 7892 2372
rect 7840 2329 7849 2363
rect 7849 2329 7883 2363
rect 7883 2329 7892 2363
rect 7840 2320 7892 2329
rect 8024 2363 8076 2372
rect 8024 2329 8033 2363
rect 8033 2329 8067 2363
rect 8067 2329 8076 2363
rect 8024 2320 8076 2329
rect 8300 2320 8352 2372
rect 4804 2252 4856 2304
rect 6552 2252 6604 2304
rect 6920 2252 6972 2304
rect 7012 2295 7064 2304
rect 7012 2261 7021 2295
rect 7021 2261 7055 2295
rect 7055 2261 7064 2295
rect 7012 2252 7064 2261
rect 7472 2252 7524 2304
rect 8116 2252 8168 2304
rect 10140 2363 10192 2372
rect 10140 2329 10149 2363
rect 10149 2329 10183 2363
rect 10183 2329 10192 2363
rect 10140 2320 10192 2329
rect 10876 2320 10928 2372
rect 14924 2388 14976 2440
rect 15476 2388 15528 2440
rect 9588 2252 9640 2304
rect 11704 2252 11756 2304
rect 13728 2295 13780 2304
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 14924 2295 14976 2304
rect 14924 2261 14933 2295
rect 14933 2261 14967 2295
rect 14967 2261 14976 2295
rect 14924 2252 14976 2261
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 16214 2150 16266 2202
rect 16278 2150 16330 2202
rect 16342 2150 16394 2202
rect 16406 2150 16458 2202
rect 16470 2150 16522 2202
rect 3700 2091 3752 2100
rect 3700 2057 3709 2091
rect 3709 2057 3743 2091
rect 3743 2057 3752 2091
rect 3700 2048 3752 2057
rect 3976 1980 4028 2032
rect 1952 1955 2004 1964
rect 1952 1921 1961 1955
rect 1961 1921 1995 1955
rect 1995 1921 2004 1955
rect 1952 1912 2004 1921
rect 3884 1912 3936 1964
rect 6736 2048 6788 2100
rect 4804 1980 4856 2032
rect 6552 1980 6604 2032
rect 9680 2048 9732 2100
rect 10876 2091 10928 2100
rect 10876 2057 10885 2091
rect 10885 2057 10919 2091
rect 10919 2057 10928 2091
rect 10876 2048 10928 2057
rect 10600 1980 10652 2032
rect 11888 1980 11940 2032
rect 14280 1980 14332 2032
rect 6368 1912 6420 1964
rect 6644 1955 6696 1964
rect 6644 1921 6653 1955
rect 6653 1921 6687 1955
rect 6687 1921 6696 1955
rect 6644 1912 6696 1921
rect 7472 1912 7524 1964
rect 8024 1912 8076 1964
rect 8392 1955 8444 1964
rect 8392 1921 8401 1955
rect 8401 1921 8435 1955
rect 8435 1921 8444 1955
rect 8392 1912 8444 1921
rect 10784 1955 10836 1964
rect 10784 1921 10793 1955
rect 10793 1921 10827 1955
rect 10827 1921 10836 1955
rect 10784 1912 10836 1921
rect 11152 1912 11204 1964
rect 11612 1912 11664 1964
rect 2596 1844 2648 1896
rect 4896 1844 4948 1896
rect 7564 1887 7616 1896
rect 4068 1708 4120 1760
rect 7564 1853 7573 1887
rect 7573 1853 7607 1887
rect 7607 1853 7616 1887
rect 7564 1844 7616 1853
rect 8668 1887 8720 1896
rect 8668 1853 8677 1887
rect 8677 1853 8711 1887
rect 8711 1853 8720 1887
rect 8668 1844 8720 1853
rect 8760 1844 8812 1896
rect 11704 1887 11756 1896
rect 5448 1776 5500 1828
rect 11704 1853 11713 1887
rect 11713 1853 11747 1887
rect 11747 1853 11756 1887
rect 11704 1844 11756 1853
rect 6552 1751 6604 1760
rect 6552 1717 6561 1751
rect 6561 1717 6595 1751
rect 6595 1717 6604 1751
rect 6552 1708 6604 1717
rect 9772 1708 9824 1760
rect 11244 1751 11296 1760
rect 11244 1717 11253 1751
rect 11253 1717 11287 1751
rect 11287 1717 11296 1751
rect 11244 1708 11296 1717
rect 13728 1887 13780 1896
rect 13728 1853 13737 1887
rect 13737 1853 13771 1887
rect 13771 1853 13780 1887
rect 13728 1844 13780 1853
rect 14556 1708 14608 1760
rect 15476 1751 15528 1760
rect 15476 1717 15485 1751
rect 15485 1717 15519 1751
rect 15519 1717 15528 1751
rect 15476 1708 15528 1717
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 1952 1504 2004 1556
rect 3884 1547 3936 1556
rect 3884 1513 3893 1547
rect 3893 1513 3927 1547
rect 3927 1513 3936 1547
rect 3884 1504 3936 1513
rect 4804 1504 4856 1556
rect 4896 1547 4948 1556
rect 4896 1513 4905 1547
rect 4905 1513 4939 1547
rect 4939 1513 4948 1547
rect 4896 1504 4948 1513
rect 6552 1504 6604 1556
rect 8116 1504 8168 1556
rect 8392 1547 8444 1556
rect 8392 1513 8401 1547
rect 8401 1513 8435 1547
rect 8435 1513 8444 1547
rect 8392 1504 8444 1513
rect 8668 1504 8720 1556
rect 9680 1504 9732 1556
rect 11244 1504 11296 1556
rect 13728 1504 13780 1556
rect 2596 1479 2648 1488
rect 2596 1445 2605 1479
rect 2605 1445 2639 1479
rect 2639 1445 2648 1479
rect 2596 1436 2648 1445
rect 10140 1436 10192 1488
rect 10600 1436 10652 1488
rect 11888 1479 11940 1488
rect 11888 1445 11897 1479
rect 11897 1445 11931 1479
rect 11931 1445 11940 1479
rect 11888 1436 11940 1445
rect 3332 1368 3384 1420
rect 6368 1368 6420 1420
rect 6736 1368 6788 1420
rect 15752 1504 15804 1556
rect 1952 1300 2004 1352
rect 2964 1343 3016 1352
rect 2964 1309 2973 1343
rect 2973 1309 3007 1343
rect 3007 1309 3016 1343
rect 2964 1300 3016 1309
rect 3700 1300 3752 1352
rect 4620 1300 4672 1352
rect 5080 1300 5132 1352
rect 5172 1232 5224 1284
rect 5448 1232 5500 1284
rect 7012 1232 7064 1284
rect 1032 1164 1084 1216
rect 6368 1164 6420 1216
rect 9496 1300 9548 1352
rect 9772 1343 9824 1352
rect 9772 1309 9781 1343
rect 9781 1309 9815 1343
rect 9815 1309 9824 1343
rect 9772 1300 9824 1309
rect 10232 1343 10284 1352
rect 10232 1309 10241 1343
rect 10241 1309 10275 1343
rect 10275 1309 10284 1343
rect 10232 1300 10284 1309
rect 9588 1232 9640 1284
rect 10784 1300 10836 1352
rect 11152 1343 11204 1352
rect 11152 1309 11161 1343
rect 11161 1309 11195 1343
rect 11195 1309 11204 1343
rect 11152 1300 11204 1309
rect 15476 1368 15528 1420
rect 12992 1232 13044 1284
rect 14924 1232 14976 1284
rect 9864 1164 9916 1216
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 16214 1062 16266 1114
rect 16278 1062 16330 1114
rect 16342 1062 16394 1114
rect 16406 1062 16458 1114
rect 16470 1062 16522 1114
<< metal2 >>
rect 1122 14362 1178 15000
rect 1122 14346 1440 14362
rect 1122 14340 1452 14346
rect 1122 14334 1400 14340
rect 1122 14200 1178 14334
rect 1400 14282 1452 14288
rect 2594 14200 2650 15000
rect 4066 14362 4122 15000
rect 3988 14334 4122 14362
rect 2134 12608 2190 12617
rect 2134 12543 2190 12552
rect 2148 12238 2176 12543
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 1504 11762 1532 12038
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 11218 1532 11698
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1320 9042 1348 9279
rect 1308 9036 1360 9042
rect 1308 8978 1360 8984
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 1228 8537 1256 8910
rect 1872 8906 1900 9386
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1214 8528 1270 8537
rect 2056 8498 2084 9862
rect 2148 8974 2176 12038
rect 2240 11558 2268 12106
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11082 2268 11494
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2240 10062 2268 11018
rect 2332 10810 2360 11018
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2608 10713 2636 14200
rect 3514 13424 3570 13433
rect 3056 13388 3108 13394
rect 3514 13359 3570 13368
rect 3056 13330 3108 13336
rect 3068 12850 3096 13330
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 2872 12368 2924 12374
rect 3148 12368 3200 12374
rect 2924 12316 3148 12322
rect 2872 12310 3200 12316
rect 2884 12294 3188 12310
rect 3252 12238 3280 12378
rect 3528 12238 3556 13359
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3620 12374 3648 12786
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3896 12306 3924 12786
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11898 3464 12038
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3700 11824 3752 11830
rect 3698 11792 3700 11801
rect 3752 11792 3754 11801
rect 3516 11756 3568 11762
rect 3698 11727 3754 11736
rect 3516 11698 3568 11704
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2594 10704 2650 10713
rect 2594 10639 2650 10648
rect 2976 10606 3004 11086
rect 3344 10674 3372 11494
rect 3528 11150 3556 11698
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3436 10810 3464 11018
rect 3896 10810 3924 12106
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 3988 10538 4016 14334
rect 4066 14200 4122 14334
rect 5538 14200 5594 15000
rect 7010 14200 7066 15000
rect 8482 14362 8538 15000
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 8482 14334 8616 14362
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 5552 13326 5580 14200
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 4080 12782 4108 13262
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12374 4660 12854
rect 4816 12714 4844 13126
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4816 12238 4844 12650
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 11150 4108 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11370 4660 11698
rect 4632 11342 4752 11370
rect 5092 11354 5120 11698
rect 4724 11286 4752 11342
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4068 11144 4120 11150
rect 4120 11104 4200 11132
rect 4068 11086 4120 11092
rect 4172 10674 4200 11104
rect 5092 10674 5120 11290
rect 5828 11150 5856 11698
rect 6564 11626 6592 12038
rect 6656 11898 6684 12174
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6564 11150 6592 11562
rect 6748 11354 6776 13262
rect 6932 12850 6960 13330
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6932 12306 6960 12786
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 6552 11144 6604 11150
rect 6828 11144 6880 11150
rect 6552 11086 6604 11092
rect 6826 11112 6828 11121
rect 6880 11112 6882 11121
rect 7024 11082 7052 14200
rect 7116 13326 7144 14282
rect 8482 14200 8538 14334
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 11898 7236 13126
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6826 11047 6882 11056
rect 7012 11076 7064 11082
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10742 5580 10950
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 1214 8463 1270 8472
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2240 8294 2268 9522
rect 3068 9178 3096 9522
rect 4632 9450 4660 9930
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3252 8974 3280 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9110 4660 9386
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4724 9042 4752 10406
rect 4816 9994 4844 10542
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10062 5580 10406
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 5552 9586 5580 9998
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5000 9178 5028 9522
rect 5828 9518 5856 9998
rect 5920 9926 5948 10610
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 5920 9722 5948 9862
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 2332 8809 2360 8910
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 2964 8832 3016 8838
rect 2318 8800 2374 8809
rect 3424 8832 3476 8838
rect 3422 8800 3424 8809
rect 3476 8800 3478 8809
rect 2964 8774 3016 8780
rect 2318 8735 2374 8744
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2240 7970 2268 8230
rect 2148 7942 2268 7970
rect 2976 7954 3004 8774
rect 3252 8758 3422 8786
rect 2964 7948 3016 7954
rect 2148 7721 2176 7942
rect 2964 7890 3016 7896
rect 3252 7886 3280 8758
rect 3422 8735 3478 8744
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 2134 7712 2190 7721
rect 2134 7647 2190 7656
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1688 6934 1716 7346
rect 1676 6928 1728 6934
rect 1676 6870 1728 6876
rect 2148 6662 2176 7346
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2240 6458 2268 7822
rect 2332 7274 2360 7822
rect 2502 7440 2558 7449
rect 2412 7404 2464 7410
rect 2502 7375 2504 7384
rect 2412 7346 2464 7352
rect 2556 7375 2558 7384
rect 2504 7346 2556 7352
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2332 6798 2360 7210
rect 2424 7002 2452 7346
rect 2608 7206 2636 7822
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2700 7410 2728 7482
rect 3238 7440 3294 7449
rect 2688 7404 2740 7410
rect 3238 7375 3240 7384
rect 2688 7346 2740 7352
rect 3292 7375 3294 7384
rect 3240 7346 3292 7352
rect 2780 7268 2832 7274
rect 2780 7210 2832 7216
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2608 6798 2636 7142
rect 2792 7002 2820 7210
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2516 6458 2544 6734
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4457 980 5170
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 938 4448 994 4457
rect 938 4383 994 4392
rect 1306 3632 1362 3641
rect 1306 3567 1362 3576
rect 1320 3534 1348 3567
rect 1688 3534 1716 4558
rect 1780 4146 1808 6258
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1872 5710 1900 6190
rect 2240 6186 2268 6258
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1872 5273 1900 5646
rect 2240 5370 2268 6122
rect 2424 5914 2452 6326
rect 2792 6089 2820 6938
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2778 6080 2834 6089
rect 2778 6015 2834 6024
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 1858 5264 1914 5273
rect 1858 5199 1914 5208
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4146 1900 4422
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1872 3602 1900 4082
rect 1964 3670 1992 4558
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4214 2820 4422
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1320 2825 1348 2926
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 1872 2446 1900 3334
rect 1964 2514 1992 3606
rect 2056 3534 2084 4082
rect 2332 3602 2360 4082
rect 2884 3738 2912 6666
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3252 6322 3280 6394
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3344 6118 3372 6258
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3344 5930 3372 6054
rect 3252 5902 3372 5930
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2976 5166 3004 5646
rect 3068 5234 3096 5646
rect 3160 5234 3188 5714
rect 3252 5370 3280 5902
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3344 5642 3372 5782
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3344 5234 3372 5578
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2976 3942 3004 5102
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2056 2650 2084 3470
rect 2332 3194 2360 3538
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2148 2854 2176 2994
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2148 2650 2176 2790
rect 2792 2650 2820 2994
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 1952 1964 2004 1970
rect 1952 1906 2004 1912
rect 1964 1562 1992 1906
rect 2596 1896 2648 1902
rect 2596 1838 2648 1844
rect 1952 1556 2004 1562
rect 1952 1498 2004 1504
rect 1964 1358 1992 1498
rect 2608 1494 2636 1838
rect 2596 1488 2648 1494
rect 2596 1430 2648 1436
rect 2976 1358 3004 2382
rect 3344 1426 3372 4626
rect 3436 4622 3464 6938
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3436 4282 3464 4558
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3436 2582 3464 2994
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3528 2009 3556 8366
rect 3620 8090 3648 8434
rect 4908 8362 4936 8842
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 4908 8022 4936 8298
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 5552 7954 5580 8774
rect 6104 8634 6132 8910
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6104 8090 6132 8570
rect 6196 8498 6224 9862
rect 6656 9674 6684 10610
rect 6564 9646 6684 9674
rect 6564 9450 6592 9646
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6196 7954 6224 8434
rect 6380 8430 6408 8842
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6472 8566 6500 8774
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6472 7954 6500 8502
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 4554 3648 6598
rect 3896 6322 3924 7754
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3974 6896 4030 6905
rect 3974 6831 4030 6840
rect 4080 6848 4108 6938
rect 4252 6860 4304 6866
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3988 6118 4016 6831
rect 4080 6820 4252 6848
rect 4252 6802 4304 6808
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4448 5710 4476 5850
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4632 5234 4660 6054
rect 4816 5914 4844 7278
rect 5000 7002 5028 7346
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 6380 6798 6408 7414
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5302 4752 5510
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4816 4758 4844 5238
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4908 4570 4936 6258
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 5370 5028 5646
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5092 5234 5120 5578
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 4528 4548 4580 4554
rect 4908 4542 5028 4570
rect 4528 4490 4580 4496
rect 4540 4146 4568 4490
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4724 4146 4752 4422
rect 4528 4140 4580 4146
rect 4712 4140 4764 4146
rect 4528 4082 4580 4088
rect 4632 4100 4712 4128
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3712 3194 3740 3402
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 4632 3058 4660 4100
rect 4712 4082 4764 4088
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4724 3194 4752 3538
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3712 2106 3740 2382
rect 3700 2100 3752 2106
rect 3700 2042 3752 2048
rect 3514 2000 3570 2009
rect 3514 1935 3570 1944
rect 3332 1420 3384 1426
rect 3332 1362 3384 1368
rect 3712 1358 3740 2042
rect 3988 2038 4016 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 3976 2032 4028 2038
rect 3976 1974 4028 1980
rect 3884 1964 3936 1970
rect 3884 1906 3936 1912
rect 3896 1562 3924 1906
rect 4080 1766 4108 2382
rect 4068 1760 4120 1766
rect 4068 1702 4120 1708
rect 4214 1660 4522 1669
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1595 4522 1604
rect 3884 1556 3936 1562
rect 3884 1498 3936 1504
rect 4632 1358 4660 2994
rect 4724 2446 4752 3130
rect 4816 3126 4844 3470
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4816 2310 4844 3062
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 4816 1562 4844 1974
rect 4896 1896 4948 1902
rect 4896 1838 4948 1844
rect 4908 1562 4936 1838
rect 4804 1556 4856 1562
rect 4804 1498 4856 1504
rect 4896 1556 4948 1562
rect 4896 1498 4948 1504
rect 1952 1352 2004 1358
rect 1952 1294 2004 1300
rect 2964 1352 3016 1358
rect 2964 1294 3016 1300
rect 3700 1352 3752 1358
rect 3700 1294 3752 1300
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 1032 1216 1084 1222
rect 1030 1184 1032 1193
rect 1084 1184 1086 1193
rect 1030 1119 1086 1128
rect 5000 800 5028 4542
rect 5092 3738 5120 5170
rect 5368 5166 5396 5782
rect 5460 5710 5488 6054
rect 6104 5778 6132 6054
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5460 5234 5488 5646
rect 6012 5370 6040 5646
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5184 4622 5212 5034
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5092 2446 5120 2926
rect 5184 2650 5212 3946
rect 5276 2854 5304 4490
rect 5368 3670 5396 5102
rect 6564 5098 6592 9386
rect 6840 9382 6868 11047
rect 7012 11018 7064 11024
rect 6918 10704 6974 10713
rect 6918 10639 6920 10648
rect 6972 10639 6974 10648
rect 6920 10610 6972 10616
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 7116 9058 7144 11086
rect 7208 9926 7236 11834
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9178 7236 9862
rect 7300 9674 7328 13194
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 11762 7512 13126
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 7760 12714 7788 12854
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7760 12374 7788 12650
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7852 12306 7880 13330
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 12850 8156 13262
rect 8214 13084 8522 13093
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13019 8522 13028
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7944 12170 7972 12310
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7944 11694 7972 12106
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11898 8064 12038
rect 8214 11996 8522 12005
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11931 8522 11940
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7654 11112 7710 11121
rect 7654 11047 7710 11056
rect 7668 10674 7696 11047
rect 7760 10674 7788 11154
rect 8036 11150 8064 11834
rect 8588 11762 8616 14334
rect 9954 14200 10010 15000
rect 11426 14200 11482 15000
rect 12898 14200 12954 15000
rect 14370 14200 14426 15000
rect 15842 14200 15898 15000
rect 17314 14200 17370 15000
rect 18786 14200 18842 15000
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8680 12986 8708 13126
rect 9140 12986 9168 13194
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9232 12782 9260 13262
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9416 12918 9444 13194
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11762 8708 12038
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8128 10810 8156 11494
rect 8496 11014 8524 11630
rect 8576 11212 8628 11218
rect 8680 11200 8708 11698
rect 8772 11354 8800 11766
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8864 11257 8892 12174
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8628 11172 8708 11200
rect 8850 11248 8906 11257
rect 8850 11183 8906 11192
rect 8576 11154 8628 11160
rect 8956 11014 8984 11630
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8214 10908 8522 10917
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10843 8522 10852
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8956 10724 8984 10950
rect 8864 10696 8984 10724
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 10130 7420 10406
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7484 9722 7512 10542
rect 7930 10432 7986 10441
rect 7930 10367 7986 10376
rect 7944 10198 7972 10367
rect 8128 10305 8156 10610
rect 8864 10606 8892 10696
rect 9048 10674 9076 11698
rect 9232 11529 9260 12174
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9218 11520 9274 11529
rect 9218 11455 9274 11464
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9140 10674 9168 11154
rect 9232 11150 9260 11455
rect 9324 11218 9352 12038
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9036 10668 9088 10674
rect 8956 10628 9036 10656
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8114 10296 8170 10305
rect 8114 10231 8170 10240
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7932 10192 7984 10198
rect 7932 10134 7984 10140
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7576 9722 7604 9930
rect 7472 9716 7524 9722
rect 7300 9646 7420 9674
rect 7472 9658 7524 9664
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7024 9030 7144 9058
rect 6918 8936 6974 8945
rect 6918 8871 6920 8880
rect 6972 8871 6974 8880
rect 6920 8842 6972 8848
rect 7024 8566 7052 9030
rect 7104 8968 7156 8974
rect 7208 8956 7236 9114
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7156 8928 7236 8956
rect 7104 8910 7156 8916
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 7116 8498 7144 8774
rect 7300 8634 7328 8978
rect 7392 8974 7420 9646
rect 7576 9568 7604 9658
rect 7484 9540 7604 9568
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7484 8430 7512 9540
rect 7668 9518 7696 10134
rect 8024 10056 8076 10062
rect 8022 10024 8024 10033
rect 8076 10024 8078 10033
rect 8022 9959 8078 9968
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7932 9580 7984 9586
rect 7984 9540 8064 9568
rect 7932 9522 7984 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 8634 7604 9386
rect 7668 8838 7696 9454
rect 7760 9024 7788 9522
rect 7932 9036 7984 9042
rect 7760 8996 7932 9024
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7478 6776 7686
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 6458 6776 6802
rect 6828 6792 6880 6798
rect 6932 6780 6960 7958
rect 7116 7954 7144 8298
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7116 7274 7144 7890
rect 7484 7750 7512 8366
rect 7576 7886 7604 8570
rect 7668 8498 7696 8774
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7760 7886 7788 8996
rect 7932 8978 7984 8984
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7852 8809 7880 8842
rect 7838 8800 7894 8809
rect 7838 8735 7894 8744
rect 8036 8566 8064 9540
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8128 8498 8156 10231
rect 8404 10062 8432 10406
rect 8392 10056 8444 10062
rect 8668 10056 8720 10062
rect 8444 10016 8616 10044
rect 8392 9998 8444 10004
rect 8214 9820 8522 9829
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9755 8522 9764
rect 8588 9518 8616 10016
rect 8668 9998 8720 10004
rect 8680 9722 8708 9998
rect 8760 9920 8812 9926
rect 8758 9888 8760 9897
rect 8812 9888 8814 9897
rect 8758 9823 8814 9832
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8864 9364 8892 10542
rect 8956 10266 8984 10628
rect 9036 10610 9088 10616
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9232 10441 9260 11086
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9218 10432 9274 10441
rect 9218 10367 9274 10376
rect 9034 10296 9090 10305
rect 8944 10260 8996 10266
rect 9324 10266 9352 10610
rect 9416 10554 9444 12038
rect 9692 11801 9720 12786
rect 9678 11792 9734 11801
rect 9678 11727 9734 11736
rect 9784 11540 9812 12786
rect 9876 12442 9904 12786
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9646 11512 9812 11540
rect 9646 11370 9674 11512
rect 9600 11342 9674 11370
rect 9600 11218 9628 11342
rect 9678 11248 9734 11257
rect 9588 11212 9640 11218
rect 9678 11183 9734 11192
rect 9588 11154 9640 11160
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9508 10674 9536 11018
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9416 10526 9628 10554
rect 9034 10231 9090 10240
rect 9312 10260 9364 10266
rect 8944 10202 8996 10208
rect 9048 10130 9076 10231
rect 9312 10202 9364 10208
rect 9416 10146 9444 10526
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9140 10118 9444 10146
rect 9140 9738 9168 10118
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9908 9260 9998
rect 9404 9920 9456 9926
rect 9232 9880 9404 9908
rect 9404 9862 9456 9868
rect 9140 9710 9352 9738
rect 9220 9648 9272 9654
rect 9218 9616 9220 9625
rect 9272 9616 9274 9625
rect 9036 9580 9088 9586
rect 9218 9551 9274 9560
rect 9036 9522 9088 9528
rect 9048 9489 9076 9522
rect 9034 9480 9090 9489
rect 9034 9415 9090 9424
rect 8944 9376 8996 9382
rect 8864 9336 8944 9364
rect 8944 9318 8996 9324
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8214 8732 8522 8741
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8667 8522 8676
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8588 8294 8616 8434
rect 8772 8401 8800 8842
rect 9324 8498 9352 9710
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9416 9586 9444 9658
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9416 9178 9444 9522
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9508 9042 9536 10202
rect 9600 10062 9628 10526
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9588 9920 9640 9926
rect 9586 9888 9588 9897
rect 9640 9888 9642 9897
rect 9586 9823 9642 9832
rect 9586 9616 9642 9625
rect 9586 9551 9588 9560
rect 9640 9551 9642 9560
rect 9588 9522 9640 9528
rect 9692 9110 9720 11183
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9784 10810 9812 11086
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9876 10742 9904 11698
rect 9968 11234 9996 14200
rect 10138 13424 10194 13433
rect 10138 13359 10194 13368
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 11898 10088 13126
rect 10152 12918 10180 13359
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10152 12073 10180 12174
rect 10138 12064 10194 12073
rect 10138 11999 10194 12008
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10060 11762 10088 11834
rect 10244 11762 10272 12786
rect 10336 12238 10364 13262
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10428 12782 10456 13194
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 12850 10640 13126
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10336 12102 10364 12174
rect 10428 12170 10456 12718
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10414 12064 10470 12073
rect 10414 11999 10470 12008
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10060 11393 10088 11698
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10046 11384 10102 11393
rect 10046 11319 10102 11328
rect 9968 11206 10088 11234
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9968 10810 9996 11086
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9770 10432 9826 10441
rect 9770 10367 9826 10376
rect 9784 10198 9812 10367
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9784 8974 9812 9930
rect 9876 9178 9904 10678
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9968 9722 9996 10610
rect 10060 10033 10088 11206
rect 10152 10538 10180 11630
rect 10244 10810 10272 11698
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10336 10577 10364 11834
rect 10428 11257 10456 11999
rect 10796 11762 10824 12106
rect 10980 11898 11008 12786
rect 11072 12306 11100 12922
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11164 12238 11192 12718
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10414 11248 10470 11257
rect 10414 11183 10470 11192
rect 10428 11150 10456 11183
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10322 10568 10378 10577
rect 10140 10532 10192 10538
rect 10428 10538 10456 11086
rect 10520 10810 10548 11698
rect 10612 11558 10640 11698
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10322 10503 10378 10512
rect 10416 10532 10468 10538
rect 10140 10474 10192 10480
rect 10416 10474 10468 10480
rect 10138 10432 10194 10441
rect 10138 10367 10194 10376
rect 10152 10062 10180 10367
rect 10232 10260 10284 10266
rect 10284 10220 10364 10248
rect 10232 10202 10284 10208
rect 10140 10056 10192 10062
rect 10046 10024 10102 10033
rect 10140 9998 10192 10004
rect 10046 9959 10102 9968
rect 10336 9761 10364 10220
rect 10428 10198 10456 10474
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10520 9994 10548 10610
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10322 9752 10378 9761
rect 9956 9716 10008 9722
rect 10322 9687 10378 9696
rect 9956 9658 10008 9664
rect 10428 9674 10456 9930
rect 10612 9926 10640 10746
rect 10704 10062 10732 11154
rect 10796 10441 10824 11698
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11257 10916 11494
rect 10874 11248 10930 11257
rect 10874 11183 10930 11192
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10980 10985 11008 11086
rect 11072 11014 11100 11086
rect 11060 11008 11112 11014
rect 10966 10976 11022 10985
rect 10888 10934 10966 10962
rect 10888 10606 10916 10934
rect 11060 10950 11112 10956
rect 10966 10911 11022 10920
rect 10876 10600 10928 10606
rect 11164 10588 11192 12038
rect 11242 11384 11298 11393
rect 11242 11319 11298 11328
rect 11256 11150 11284 11319
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11348 10742 11376 10950
rect 11336 10736 11388 10742
rect 11440 10713 11468 14200
rect 12214 13628 12522 13637
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13563 12522 13572
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12176 12918 12204 13126
rect 12268 12986 12296 13466
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12728 12782 12756 13262
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12214 12540 12522 12549
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12475 12522 12484
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 11532 11762 11560 12174
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11336 10678 11388 10684
rect 11426 10704 11482 10713
rect 11426 10639 11482 10648
rect 10876 10542 10928 10548
rect 11072 10560 11192 10588
rect 10782 10432 10838 10441
rect 10782 10367 10838 10376
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10428 9654 10732 9674
rect 10428 9648 10744 9654
rect 10428 9646 10692 9648
rect 9954 9616 10010 9625
rect 10692 9590 10744 9596
rect 9954 9551 10010 9560
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9678 8664 9734 8673
rect 9678 8599 9734 8608
rect 9586 8528 9642 8537
rect 9312 8492 9364 8498
rect 9692 8498 9720 8599
rect 9772 8560 9824 8566
rect 9876 8548 9904 9114
rect 9968 8974 9996 9551
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10152 8974 10180 9386
rect 10704 8974 10732 9590
rect 10888 9489 10916 9862
rect 11072 9674 11100 10560
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 10305 11192 10406
rect 11150 10296 11206 10305
rect 11150 10231 11206 10240
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11440 10062 11468 10134
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 10980 9646 11100 9674
rect 10874 9480 10930 9489
rect 10874 9415 10930 9424
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 9954 8800 10010 8809
rect 9954 8735 10010 8744
rect 9824 8520 9904 8548
rect 9772 8502 9824 8508
rect 9586 8463 9588 8472
rect 9312 8434 9364 8440
rect 9640 8463 9642 8472
rect 9680 8492 9732 8498
rect 9588 8434 9640 8440
rect 9680 8434 9732 8440
rect 8758 8392 8814 8401
rect 8758 8327 8814 8336
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8036 7954 8340 7970
rect 8024 7948 8352 7954
rect 8076 7942 8300 7948
rect 8024 7890 8076 7896
rect 8300 7890 8352 7896
rect 8404 7886 8432 8230
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7410 7880 7686
rect 8128 7546 8156 7822
rect 8214 7644 8522 7653
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7579 8522 7588
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8588 7410 8616 8230
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7024 6934 7052 7142
rect 8128 6934 8156 7346
rect 8772 7274 8800 8327
rect 9324 8022 9352 8434
rect 9864 8424 9916 8430
rect 9784 8384 9864 8412
rect 9496 8356 9548 8362
rect 9784 8312 9812 8384
rect 9864 8366 9916 8372
rect 9496 8298 9548 8304
rect 9772 8306 9824 8312
rect 9508 8090 9536 8298
rect 9772 8248 9824 8254
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9324 7410 9352 7958
rect 9968 7954 9996 8735
rect 10244 8566 10272 8842
rect 10692 8832 10744 8838
rect 10796 8809 10824 8842
rect 10692 8774 10744 8780
rect 10782 8800 10838 8809
rect 10232 8560 10284 8566
rect 10138 8528 10194 8537
rect 10048 8492 10100 8498
rect 10232 8502 10284 8508
rect 10322 8528 10378 8537
rect 10138 8463 10194 8472
rect 10704 8498 10732 8774
rect 10782 8735 10838 8744
rect 10322 8463 10378 8472
rect 10508 8492 10560 8498
rect 10048 8434 10100 8440
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 6880 6752 6960 6780
rect 6828 6734 6880 6740
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 5166 6684 6258
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6748 5234 6776 6122
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7116 5778 7144 6054
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4690 6500 4966
rect 6656 4826 6684 5102
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5644 4214 5672 4558
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 5920 3194 5948 3470
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 5092 1358 5120 2382
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 5172 1284 5224 1290
rect 5276 1272 5304 2790
rect 5460 2428 5488 2994
rect 5920 2446 5948 3130
rect 6012 2650 6040 3470
rect 6380 2650 6408 4014
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 5540 2440 5592 2446
rect 5460 2400 5540 2428
rect 5460 1834 5488 2400
rect 5540 2382 5592 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6564 2038 6592 2246
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6656 1970 6684 4626
rect 6748 3398 6776 5170
rect 6840 4214 6868 5646
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7012 5160 7064 5166
rect 6932 5120 7012 5148
rect 6932 4690 6960 5120
rect 7012 5102 7064 5108
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6920 4480 6972 4486
rect 7024 4468 7052 4694
rect 6972 4440 7052 4468
rect 6920 4422 6972 4428
rect 6828 4208 6880 4214
rect 6880 4156 6960 4162
rect 6828 4150 6960 4156
rect 6840 4134 6960 4150
rect 7024 4146 7052 4440
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6736 3120 6788 3126
rect 6840 3108 6868 3470
rect 6788 3080 6868 3108
rect 6736 3062 6788 3068
rect 6932 2774 6960 4134
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7024 2938 7052 4082
rect 7116 4078 7144 5102
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7576 4486 7604 4762
rect 7944 4622 7972 5170
rect 8036 4672 8064 6598
rect 8128 6254 8156 6870
rect 8496 6798 8524 7142
rect 9600 6866 9628 7414
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8214 6556 8522 6565
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6491 8522 6500
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8588 5914 8616 6258
rect 8772 6186 8800 6666
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8128 5370 8156 5578
rect 8214 5468 8522 5477
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5403 8522 5412
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8036 4644 8156 4672
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7576 4214 7604 4422
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 8128 4078 8156 4644
rect 8220 4622 8248 5102
rect 8680 4690 8708 6054
rect 8772 5234 8800 6122
rect 8864 5370 8892 6258
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8956 5166 8984 5510
rect 9140 5302 9168 5646
rect 9324 5302 9352 6598
rect 9600 6186 9628 6802
rect 9692 6662 9720 7686
rect 10060 7342 10088 8434
rect 10152 8362 10180 8463
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10336 8294 10364 8463
rect 10508 8434 10560 8440
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10244 8266 10364 8294
rect 10416 8288 10468 8294
rect 10244 7886 10272 8266
rect 10416 8230 10468 8236
rect 10428 7954 10456 8230
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 10060 6390 10088 6666
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10152 6322 10180 7822
rect 10244 7546 10272 7822
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10428 7478 10456 7890
rect 10520 7818 10548 8434
rect 10704 8362 10732 8434
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10520 6458 10548 7754
rect 10796 6458 10824 8434
rect 10888 6934 10916 8978
rect 10980 8838 11008 9646
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 11440 8498 11468 9998
rect 11532 9926 11560 11698
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 11076 11664 11082
rect 11716 11064 11744 11290
rect 11808 11150 11836 12106
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11796 11144 11848 11150
rect 11664 11036 11744 11064
rect 11794 11112 11796 11121
rect 11848 11112 11850 11121
rect 11794 11047 11850 11056
rect 11612 11018 11664 11024
rect 11808 11014 11836 11047
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11900 10713 11928 11766
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11992 11257 12020 11630
rect 11978 11248 12034 11257
rect 11978 11183 12034 11192
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11886 10704 11942 10713
rect 11612 10668 11664 10674
rect 11886 10639 11942 10648
rect 11612 10610 11664 10616
rect 11624 9926 11652 10610
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11900 10441 11928 10542
rect 11886 10432 11942 10441
rect 11886 10367 11942 10376
rect 11900 10266 11928 10367
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11992 10112 12020 10746
rect 12084 10674 12112 11698
rect 12544 11665 12572 11698
rect 12530 11656 12586 11665
rect 12530 11591 12586 11600
rect 12214 11452 12522 11461
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11387 12522 11396
rect 12636 11354 12664 12174
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12636 11218 12664 11290
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12440 11144 12492 11150
rect 12492 11104 12572 11132
rect 12440 11086 12492 11092
rect 12544 11098 12572 11104
rect 12728 11098 12756 12038
rect 12912 11762 12940 14200
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 12986 13400 13126
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13188 12442 13216 12922
rect 13464 12866 13492 13262
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13372 12838 13492 12866
rect 13372 12782 13400 12838
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13372 12442 13400 12718
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 12990 11792 13046 11801
rect 12900 11756 12952 11762
rect 12990 11727 12992 11736
rect 12900 11698 12952 11704
rect 13044 11727 13046 11736
rect 12992 11698 13044 11704
rect 12806 11656 12862 11665
rect 12806 11591 12862 11600
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11900 10084 12020 10112
rect 11796 10056 11848 10062
rect 11900 10044 11928 10084
rect 11848 10016 11928 10044
rect 11796 9998 11848 10004
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11612 9920 11664 9926
rect 11900 9897 11928 10016
rect 11612 9862 11664 9868
rect 11886 9888 11942 9897
rect 11624 9625 11652 9862
rect 11886 9823 11942 9832
rect 11978 9752 12034 9761
rect 12084 9722 12112 10610
rect 12268 10470 12296 11086
rect 12544 11070 12756 11098
rect 12544 10606 12572 11070
rect 12820 10810 12848 11591
rect 13096 11218 13124 12378
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12214 10364 12522 10373
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10299 12522 10308
rect 12636 10266 12664 10474
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10266 12756 10406
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12820 10146 12848 10610
rect 12912 10282 12940 10950
rect 13188 10674 13216 11290
rect 13372 11257 13400 11290
rect 13358 11248 13414 11257
rect 13358 11183 13414 11192
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13280 10538 13308 10950
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 12912 10254 13032 10282
rect 12624 10124 12676 10130
rect 12820 10118 12940 10146
rect 12624 10066 12676 10072
rect 11978 9687 12034 9696
rect 12072 9716 12124 9722
rect 11610 9616 11666 9625
rect 11992 9586 12020 9687
rect 12072 9658 12124 9664
rect 12636 9586 12664 10066
rect 12912 10062 12940 10118
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 11610 9551 11666 9560
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 7546 11008 8298
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10980 6866 11008 7482
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11072 6798 11100 8434
rect 11624 8401 11652 9318
rect 11716 9178 11744 9522
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11716 8974 11744 9114
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11900 8430 11928 9386
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11888 8424 11940 8430
rect 11610 8392 11666 8401
rect 11992 8401 12020 8842
rect 12084 8809 12112 9454
rect 12214 9276 12522 9285
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9211 12522 9220
rect 12530 9072 12586 9081
rect 12530 9007 12532 9016
rect 12584 9007 12586 9016
rect 12532 8978 12584 8984
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8809 12664 8910
rect 12070 8800 12126 8809
rect 12070 8735 12126 8744
rect 12622 8800 12678 8809
rect 12622 8735 12678 8744
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 11888 8366 11940 8372
rect 11978 8392 12034 8401
rect 11610 8327 11666 8336
rect 11624 8294 11652 8327
rect 11624 8288 11848 8294
rect 11624 8266 11796 8288
rect 11796 8230 11848 8236
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11256 7857 11284 8026
rect 11808 7886 11836 8230
rect 11796 7880 11848 7886
rect 11242 7848 11298 7857
rect 11796 7822 11848 7828
rect 11242 7783 11298 7792
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6662 11100 6734
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9600 5914 9628 6122
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9876 5710 9904 6258
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10336 5710 10364 6122
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9692 5302 9720 5510
rect 9876 5370 9904 5646
rect 11072 5370 11100 6598
rect 11256 6322 11284 7783
rect 11900 7410 11928 8366
rect 12084 8362 12112 8502
rect 12728 8498 12756 9590
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 11978 8327 12034 8336
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12084 7954 12112 8298
rect 12214 8188 12522 8197
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8123 12522 8132
rect 12728 8090 12756 8434
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12820 7818 12848 9930
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12912 8974 12940 9658
rect 13004 9586 13032 10254
rect 13096 10198 13124 10474
rect 13084 10192 13136 10198
rect 13372 10146 13400 10610
rect 13084 10134 13136 10140
rect 13280 10118 13400 10146
rect 13280 10062 13308 10118
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9654 13124 9862
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13004 9178 13032 9522
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12912 8022 12940 8910
rect 13084 8832 13136 8838
rect 13004 8780 13084 8786
rect 13004 8774 13136 8780
rect 13004 8758 13124 8774
rect 13004 8498 13032 8758
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5710 11836 6054
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8956 4826 8984 5102
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8956 4622 8984 4762
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 9784 4554 9812 4966
rect 9876 4826 9904 5306
rect 11624 5234 11652 5578
rect 11900 5302 11928 7210
rect 12084 6730 12112 7346
rect 12214 7100 12522 7109
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7035 12522 7044
rect 12728 6798 12756 7686
rect 13004 7342 13032 8434
rect 13188 7936 13216 9998
rect 13280 9568 13308 9998
rect 13360 9580 13412 9586
rect 13280 9540 13360 9568
rect 13360 9522 13412 9528
rect 13266 9480 13322 9489
rect 13372 9450 13400 9522
rect 13464 9450 13492 11766
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 10985 13584 11494
rect 13648 11082 13676 13126
rect 14384 12918 14412 14200
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14476 12850 14504 13262
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14108 12238 14136 12718
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14002 11928 14058 11937
rect 14002 11863 14058 11872
rect 14016 11694 14044 11863
rect 14200 11762 14228 12174
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13542 10976 13598 10985
rect 13542 10911 13598 10920
rect 13556 10674 13584 10911
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13648 9586 13676 10542
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 9722 13768 10406
rect 13832 10062 13860 11562
rect 14384 11558 14412 12106
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13924 9926 13952 10610
rect 14186 10160 14242 10169
rect 14186 10095 14242 10104
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 14108 9654 14136 9930
rect 14200 9654 14228 10095
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13266 9415 13322 9424
rect 13360 9444 13412 9450
rect 13280 8974 13308 9415
rect 13360 9386 13412 9392
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13372 8838 13400 9386
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13280 8294 13308 8570
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13096 7908 13216 7936
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13096 7018 13124 7908
rect 13280 7886 13308 8230
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13004 6990 13124 7018
rect 12716 6792 12768 6798
rect 12636 6752 12716 6780
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 12214 6012 12522 6021
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5947 12522 5956
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11624 4826 11652 5170
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 8214 4380 8522 4389
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4315 8522 4324
rect 11164 4282 11192 4762
rect 11992 4706 12020 5714
rect 12636 5710 12664 6752
rect 12716 6734 12768 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 6322 12848 6598
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12728 5914 12756 6258
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12912 5710 12940 6734
rect 13004 6118 13032 6990
rect 13084 6928 13136 6934
rect 13084 6870 13136 6876
rect 13096 6322 13124 6870
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12214 4924 12522 4933
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4859 12522 4868
rect 12636 4826 12664 5238
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 11900 4678 12020 4706
rect 12440 4684 12492 4690
rect 11900 4622 11928 4678
rect 12440 4626 12492 4632
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 7104 4072 7156 4078
rect 7472 4072 7524 4078
rect 7156 4032 7236 4060
rect 7104 4014 7156 4020
rect 7024 2910 7144 2938
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6748 2746 6960 2774
rect 6748 2106 6776 2746
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6932 2310 6960 2586
rect 7024 2446 7052 2790
rect 7116 2446 7144 2910
rect 7208 2854 7236 4032
rect 7472 4014 7524 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 7484 3738 7512 4014
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8036 3738 8064 3878
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8128 3602 8156 4014
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7760 3194 7788 3470
rect 8214 3292 8522 3301
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3227 8522 3236
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7484 2514 7512 2790
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 6368 1964 6420 1970
rect 6368 1906 6420 1912
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 5448 1828 5500 1834
rect 5448 1770 5500 1776
rect 5460 1290 5488 1770
rect 6380 1426 6408 1906
rect 6552 1760 6604 1766
rect 6552 1702 6604 1708
rect 6564 1562 6592 1702
rect 6552 1556 6604 1562
rect 6552 1498 6604 1504
rect 6748 1426 6776 2042
rect 6368 1420 6420 1426
rect 6368 1362 6420 1368
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 5224 1244 5304 1272
rect 5448 1284 5500 1290
rect 5172 1226 5224 1232
rect 5448 1226 5500 1232
rect 6380 1222 6408 1362
rect 7024 1290 7052 2246
rect 7484 1970 7512 2246
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7576 1902 7604 2382
rect 7852 2378 7880 3062
rect 8496 2922 8524 3062
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8036 2378 8064 2450
rect 8312 2378 8340 2790
rect 8680 2446 8708 3062
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8036 1970 8064 2314
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8024 1964 8076 1970
rect 8024 1906 8076 1912
rect 7564 1896 7616 1902
rect 7564 1838 7616 1844
rect 8128 1562 8156 2246
rect 8214 2204 8522 2213
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2139 8522 2148
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 8404 1562 8432 1906
rect 8772 1902 8800 2790
rect 9048 2446 9076 3130
rect 9232 3058 9260 4014
rect 9416 3602 9444 4014
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8668 1896 8720 1902
rect 8668 1838 8720 1844
rect 8760 1896 8812 1902
rect 8760 1838 8812 1844
rect 8680 1562 8708 1838
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 8392 1556 8444 1562
rect 8392 1498 8444 1504
rect 8668 1556 8720 1562
rect 8668 1498 8720 1504
rect 9508 1358 9536 3606
rect 9600 3534 9628 4082
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9784 3942 9812 4014
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9600 3194 9628 3470
rect 9692 3194 9720 3470
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9784 3058 9812 3878
rect 9968 3670 9996 3878
rect 10152 3738 10180 4082
rect 11164 4010 11192 4218
rect 11900 4146 11928 4558
rect 12452 4486 12480 4626
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 11888 4140 11940 4146
rect 11624 4100 11888 4128
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10152 3618 10180 3674
rect 9968 3534 9996 3606
rect 10152 3590 10272 3618
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 9600 1290 9628 2246
rect 9692 2106 9720 2382
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9692 1562 9720 2042
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 9680 1556 9732 1562
rect 9680 1498 9732 1504
rect 9784 1358 9812 1702
rect 9772 1352 9824 1358
rect 9772 1294 9824 1300
rect 7012 1284 7064 1290
rect 7012 1226 7064 1232
rect 9588 1284 9640 1290
rect 9588 1226 9640 1232
rect 9876 1222 9904 2586
rect 10152 2514 10180 3470
rect 10244 2990 10272 3590
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10796 2650 10824 3878
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11152 2984 11204 2990
rect 10980 2932 11152 2938
rect 10980 2926 11204 2932
rect 10980 2922 11192 2926
rect 10968 2916 11192 2922
rect 11020 2910 11192 2916
rect 10968 2858 11020 2864
rect 11256 2650 11284 2994
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 10152 1494 10180 2314
rect 10140 1488 10192 1494
rect 10140 1430 10192 1436
rect 10244 1358 10272 2450
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10888 2106 10916 2314
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10600 2032 10652 2038
rect 10600 1974 10652 1980
rect 10612 1494 10640 1974
rect 11624 1970 11652 4100
rect 11888 4082 11940 4088
rect 12452 4078 12480 4422
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3466 11836 3878
rect 12084 3738 12112 3946
rect 12214 3836 12522 3845
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3771 12522 3780
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 12084 3126 12112 3674
rect 13004 3398 13032 6054
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13096 5166 13124 5646
rect 13188 5370 13216 7754
rect 13372 7546 13400 8434
rect 13464 8362 13492 8910
rect 13556 8566 13584 9522
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13648 9110 13676 9386
rect 13636 9104 13688 9110
rect 14292 9092 14320 10610
rect 14476 9654 14504 12786
rect 14568 12782 14596 13194
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14752 12442 14780 13194
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15304 12850 15332 13126
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11898 14596 12038
rect 14844 11898 14872 12174
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 15212 11762 15240 12786
rect 15488 12646 15516 12922
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12238 15516 12582
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15212 11150 15240 11494
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 14752 10810 14780 11086
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 15212 10742 15240 10950
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 14844 9994 14872 10678
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14200 9081 14320 9092
rect 13636 9046 13688 9052
rect 14186 9072 14320 9081
rect 14242 9064 14320 9072
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14186 9007 14242 9016
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 14200 8498 14228 9007
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13464 7410 13492 7822
rect 13740 7478 13768 7822
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13832 7342 13860 8298
rect 13924 8294 13952 8434
rect 14292 8362 14320 8774
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7954 13952 8230
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 14384 7886 14412 8570
rect 14476 8537 14504 9046
rect 14568 9042 14596 9658
rect 14844 9110 14872 9930
rect 14936 9450 14964 10542
rect 15028 10198 15056 10610
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15016 10192 15068 10198
rect 15016 10134 15068 10140
rect 15014 9888 15070 9897
rect 15212 9874 15240 10542
rect 15304 10266 15332 11154
rect 15488 10742 15516 11222
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15396 10441 15424 10678
rect 15580 10588 15608 11494
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15672 10810 15700 10950
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15488 10560 15608 10588
rect 15382 10432 15438 10441
rect 15382 10367 15438 10376
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15070 9846 15240 9874
rect 15014 9823 15070 9832
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14936 8974 14964 9386
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14554 8800 14610 8809
rect 14554 8735 14610 8744
rect 14568 8634 14596 8735
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14462 8528 14518 8537
rect 14462 8463 14464 8472
rect 14516 8463 14518 8472
rect 14464 8434 14516 8440
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13280 6390 13308 7278
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14292 6866 14320 7210
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13372 6254 13400 6734
rect 14568 6662 14596 8570
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14660 7886 14688 8230
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13372 5710 13400 5850
rect 13924 5778 13952 6054
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13924 5302 13952 5714
rect 14016 5302 14044 6122
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14108 5302 14136 5578
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13096 4826 13124 5102
rect 13924 4826 13952 5238
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13924 4282 13952 4762
rect 14384 4554 14412 6054
rect 14476 5778 14504 6598
rect 14568 5778 14596 6598
rect 14660 6390 14688 6598
rect 14752 6458 14780 7890
rect 15028 7886 15056 9823
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15120 7274 15148 9522
rect 15212 8634 15240 9522
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15198 8392 15254 8401
rect 15198 8327 15254 8336
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14844 6254 14872 6802
rect 15120 6390 15148 7210
rect 15212 6798 15240 8327
rect 15304 7410 15332 9658
rect 15488 9654 15516 10560
rect 15566 10160 15622 10169
rect 15566 10095 15622 10104
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15384 9172 15436 9178
rect 15488 9160 15516 9590
rect 15436 9132 15516 9160
rect 15384 9114 15436 9120
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 15212 4826 15240 6734
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13096 3534 13124 4014
rect 13924 3602 13952 4218
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12992 3120 13044 3126
rect 12992 3062 13044 3068
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11716 2310 11744 2994
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 2854 12112 2926
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12214 2748 12522 2757
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2683 12522 2692
rect 13004 2650 13032 3062
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13096 2530 13124 3470
rect 13924 3194 13952 3538
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13004 2502 13124 2530
rect 13004 2446 13032 2502
rect 14936 2446 14964 3674
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11612 1964 11664 1970
rect 11612 1906 11664 1912
rect 10600 1488 10652 1494
rect 10600 1430 10652 1436
rect 10796 1358 10824 1906
rect 11164 1358 11192 1906
rect 11716 1902 11744 2246
rect 11888 2032 11940 2038
rect 11888 1974 11940 1980
rect 11704 1896 11756 1902
rect 11704 1838 11756 1844
rect 11244 1760 11296 1766
rect 11244 1702 11296 1708
rect 11256 1562 11284 1702
rect 11244 1556 11296 1562
rect 11244 1498 11296 1504
rect 11900 1494 11928 1974
rect 12214 1660 12522 1669
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1595 12522 1604
rect 11888 1488 11940 1494
rect 11888 1430 11940 1436
rect 10232 1352 10284 1358
rect 10232 1294 10284 1300
rect 10784 1352 10836 1358
rect 10784 1294 10836 1300
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 13004 1290 13032 2382
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 13740 1902 13768 2246
rect 14292 2038 14320 2246
rect 14280 2032 14332 2038
rect 14280 1974 14332 1980
rect 13728 1896 13780 1902
rect 13728 1838 13780 1844
rect 13740 1562 13768 1838
rect 14556 1760 14608 1766
rect 14556 1702 14608 1708
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 12992 1284 13044 1290
rect 12992 1226 13044 1232
rect 6368 1216 6420 1222
rect 6368 1158 6420 1164
rect 9864 1216 9916 1222
rect 9864 1158 9916 1164
rect 8214 1116 8522 1125
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1051 8522 1060
rect 4986 0 5042 800
rect 14568 762 14596 1702
rect 14936 1290 14964 2246
rect 15396 1329 15424 8910
rect 15488 8498 15516 8910
rect 15580 8537 15608 10095
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15566 8528 15622 8537
rect 15476 8492 15528 8498
rect 15566 8463 15622 8472
rect 15476 8434 15528 8440
rect 15566 8392 15622 8401
rect 15672 8378 15700 9998
rect 15764 9450 15792 11086
rect 15856 11082 15884 14200
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15948 11558 15976 12786
rect 16132 12782 16160 13194
rect 16214 13084 16522 13093
rect 16214 13082 16220 13084
rect 16276 13082 16300 13084
rect 16356 13082 16380 13084
rect 16436 13082 16460 13084
rect 16516 13082 16522 13084
rect 16276 13030 16278 13082
rect 16458 13030 16460 13082
rect 16214 13028 16220 13030
rect 16276 13028 16300 13030
rect 16356 13028 16380 13030
rect 16436 13028 16460 13030
rect 16516 13028 16522 13030
rect 16214 13019 16522 13028
rect 16684 12918 16712 13262
rect 16776 12986 16804 13262
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 12238 16160 12718
rect 16776 12238 16804 12786
rect 17328 12434 17356 14200
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17420 12442 17448 13194
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17052 12406 17356 12434
rect 17408 12436 17460 12442
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16214 11996 16522 12005
rect 16214 11994 16220 11996
rect 16276 11994 16300 11996
rect 16356 11994 16380 11996
rect 16436 11994 16460 11996
rect 16516 11994 16522 11996
rect 16276 11942 16278 11994
rect 16458 11942 16460 11994
rect 16214 11940 16220 11942
rect 16276 11940 16300 11942
rect 16356 11940 16380 11942
rect 16436 11940 16460 11942
rect 16516 11940 16522 11942
rect 16214 11931 16522 11940
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11286 16252 11494
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10606 15976 10950
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15622 8350 15700 8378
rect 15566 8327 15622 8336
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15488 7478 15516 7958
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15488 5370 15516 6666
rect 15580 6662 15608 8327
rect 15764 8022 15792 8842
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15856 8634 15884 8774
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15948 8514 15976 9386
rect 15856 8486 15976 8514
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 6798 15792 7142
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6322 15792 6598
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15856 6089 15884 8486
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15948 7478 15976 8230
rect 16040 7954 16068 11222
rect 16304 11144 16356 11150
rect 16302 11112 16304 11121
rect 16356 11112 16358 11121
rect 16120 11076 16172 11082
rect 16302 11047 16358 11056
rect 16120 11018 16172 11024
rect 16132 10538 16160 11018
rect 16214 10908 16522 10917
rect 16214 10906 16220 10908
rect 16276 10906 16300 10908
rect 16356 10906 16380 10908
rect 16436 10906 16460 10908
rect 16516 10906 16522 10908
rect 16276 10854 16278 10906
rect 16458 10854 16460 10906
rect 16214 10852 16220 10854
rect 16276 10852 16300 10854
rect 16356 10852 16380 10854
rect 16436 10852 16460 10854
rect 16516 10852 16522 10854
rect 16214 10843 16522 10852
rect 16854 10704 16910 10713
rect 16854 10639 16910 10648
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16776 10062 16804 10542
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16214 9820 16522 9829
rect 16214 9818 16220 9820
rect 16276 9818 16300 9820
rect 16356 9818 16380 9820
rect 16436 9818 16460 9820
rect 16516 9818 16522 9820
rect 16276 9766 16278 9818
rect 16458 9766 16460 9818
rect 16214 9764 16220 9766
rect 16276 9764 16300 9766
rect 16356 9764 16380 9766
rect 16436 9764 16460 9766
rect 16516 9764 16522 9766
rect 16214 9755 16522 9764
rect 16776 9654 16804 9998
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16214 8732 16522 8741
rect 16214 8730 16220 8732
rect 16276 8730 16300 8732
rect 16356 8730 16380 8732
rect 16436 8730 16460 8732
rect 16516 8730 16522 8732
rect 16276 8678 16278 8730
rect 16458 8678 16460 8730
rect 16214 8676 16220 8678
rect 16276 8676 16300 8678
rect 16356 8676 16380 8678
rect 16436 8676 16460 8678
rect 16516 8676 16522 8678
rect 16214 8667 16522 8676
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 15948 6474 15976 7414
rect 16040 7410 16068 7890
rect 16592 7886 16620 8230
rect 16580 7880 16632 7886
rect 16210 7848 16266 7857
rect 16580 7822 16632 7828
rect 16132 7792 16210 7800
rect 16132 7772 16212 7792
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16132 6798 16160 7772
rect 16264 7783 16266 7792
rect 16212 7754 16264 7760
rect 16214 7644 16522 7653
rect 16214 7642 16220 7644
rect 16276 7642 16300 7644
rect 16356 7642 16380 7644
rect 16436 7642 16460 7644
rect 16516 7642 16522 7644
rect 16276 7590 16278 7642
rect 16458 7590 16460 7642
rect 16214 7588 16220 7590
rect 16276 7588 16300 7590
rect 16356 7588 16380 7590
rect 16436 7588 16460 7590
rect 16516 7588 16522 7590
rect 16214 7579 16522 7588
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16214 6556 16522 6565
rect 16214 6554 16220 6556
rect 16276 6554 16300 6556
rect 16356 6554 16380 6556
rect 16436 6554 16460 6556
rect 16516 6554 16522 6556
rect 16276 6502 16278 6554
rect 16458 6502 16460 6554
rect 16214 6500 16220 6502
rect 16276 6500 16300 6502
rect 16356 6500 16380 6502
rect 16436 6500 16460 6502
rect 16516 6500 16522 6502
rect 16214 6491 16522 6500
rect 15948 6446 16160 6474
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15842 6080 15898 6089
rect 15842 6015 15898 6024
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15856 4146 15884 5170
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15856 3058 15884 4082
rect 15948 3641 15976 6122
rect 16040 5914 16068 6258
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16040 5250 16068 5850
rect 16132 5778 16160 6446
rect 16592 5778 16620 6734
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16132 5370 16160 5714
rect 16214 5468 16522 5477
rect 16214 5466 16220 5468
rect 16276 5466 16300 5468
rect 16356 5466 16380 5468
rect 16436 5466 16460 5468
rect 16516 5466 16522 5468
rect 16276 5414 16278 5466
rect 16458 5414 16460 5466
rect 16214 5412 16220 5414
rect 16276 5412 16300 5414
rect 16356 5412 16380 5414
rect 16436 5412 16460 5414
rect 16516 5412 16522 5414
rect 16214 5403 16522 5412
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16040 5234 16160 5250
rect 16684 5234 16712 8366
rect 16776 7546 16804 8910
rect 16868 7886 16896 10639
rect 17052 10130 17080 12406
rect 17408 12378 17460 12384
rect 17420 12238 17448 12378
rect 17604 12306 17632 13126
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17696 12442 17724 12854
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17236 10674 17264 11698
rect 17328 11354 17356 12174
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11762 17448 12038
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17420 11150 17448 11698
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 18064 11082 18092 12786
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17144 8974 17172 9522
rect 17236 9178 17264 10474
rect 17972 10198 18000 10746
rect 18156 10742 18184 11494
rect 18248 10742 18276 12582
rect 18800 12374 18828 14200
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17420 9586 17448 9930
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17420 9042 17448 9522
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 9110 17632 9318
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17132 8968 17184 8974
rect 17130 8936 17132 8945
rect 17184 8936 17186 8945
rect 17130 8871 17186 8880
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16868 7342 16896 7822
rect 16960 7818 16988 8570
rect 17604 8566 17632 9046
rect 17972 8974 18000 10134
rect 18156 10062 18184 10678
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17788 7886 17816 8298
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16960 7410 16988 7754
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16856 6792 16908 6798
rect 16960 6780 16988 7346
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16908 6752 16988 6780
rect 16856 6734 16908 6740
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 16868 5370 16896 5578
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16040 5228 16172 5234
rect 16040 5222 16120 5228
rect 16120 5170 16172 5176
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16040 4554 16068 4966
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 16214 4380 16522 4389
rect 16214 4378 16220 4380
rect 16276 4378 16300 4380
rect 16356 4378 16380 4380
rect 16436 4378 16460 4380
rect 16516 4378 16522 4380
rect 16276 4326 16278 4378
rect 16458 4326 16460 4378
rect 16214 4324 16220 4326
rect 16276 4324 16300 4326
rect 16356 4324 16380 4326
rect 16436 4324 16460 4326
rect 16516 4324 16522 4326
rect 16214 4315 16522 4324
rect 16960 4146 16988 5170
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16592 3738 16620 4082
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 15934 3632 15990 3641
rect 15934 3567 15990 3576
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15580 2514 15608 2994
rect 16040 2854 16068 3470
rect 16214 3292 16522 3301
rect 16214 3290 16220 3292
rect 16276 3290 16300 3292
rect 16356 3290 16380 3292
rect 16436 3290 16460 3292
rect 16516 3290 16522 3292
rect 16276 3238 16278 3290
rect 16458 3238 16460 3290
rect 16214 3236 16220 3238
rect 16276 3236 16300 3238
rect 16356 3236 16380 3238
rect 16436 3236 16460 3238
rect 16516 3236 16522 3238
rect 16214 3227 16522 3236
rect 16592 3058 16620 3674
rect 16684 3534 16712 3878
rect 17052 3738 17080 6938
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17328 6458 17356 6734
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17328 6322 17356 6394
rect 17788 6390 17816 7822
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18156 7410 18184 7686
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18340 6662 18368 7822
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17788 5710 17816 6326
rect 18340 6186 18368 6598
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18432 5914 18460 6734
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17236 5370 17264 5646
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17144 3534 17172 4082
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17420 3602 17448 4014
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 3194 16712 3334
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 17420 3058 17448 3538
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 17696 2582 17724 2994
rect 17684 2576 17736 2582
rect 17684 2518 17736 2524
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15488 1766 15516 2382
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 15488 1426 15516 1702
rect 15764 1562 15792 2450
rect 16214 2204 16522 2213
rect 16214 2202 16220 2204
rect 16276 2202 16300 2204
rect 16356 2202 16380 2204
rect 16436 2202 16460 2204
rect 16516 2202 16522 2204
rect 16276 2150 16278 2202
rect 16458 2150 16460 2202
rect 16214 2148 16220 2150
rect 16276 2148 16300 2150
rect 16356 2148 16380 2150
rect 16436 2148 16460 2150
rect 16516 2148 16522 2150
rect 16214 2139 16522 2148
rect 15752 1556 15804 1562
rect 15752 1498 15804 1504
rect 15476 1420 15528 1426
rect 15476 1362 15528 1368
rect 15382 1320 15438 1329
rect 14924 1284 14976 1290
rect 15382 1255 15438 1264
rect 14924 1226 14976 1232
rect 16214 1116 16522 1125
rect 16214 1114 16220 1116
rect 16276 1114 16300 1116
rect 16356 1114 16380 1116
rect 16436 1114 16460 1116
rect 16516 1114 16522 1116
rect 16276 1062 16278 1114
rect 16458 1062 16460 1114
rect 16214 1060 16220 1062
rect 16276 1060 16300 1062
rect 16356 1060 16380 1062
rect 16436 1060 16460 1062
rect 16516 1060 16522 1062
rect 16214 1051 16522 1060
rect 14844 870 14964 898
rect 14844 762 14872 870
rect 14936 800 14964 870
rect 14568 734 14872 762
rect 14922 0 14978 800
<< via2 >>
rect 2134 12552 2190 12608
rect 1306 9288 1362 9344
rect 1214 8472 1270 8528
rect 3514 13368 3570 13424
rect 3698 11772 3700 11792
rect 3700 11772 3752 11792
rect 3752 11772 3754 11792
rect 3698 11736 3754 11772
rect 2594 10648 2650 10704
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 6826 11092 6828 11112
rect 6828 11092 6880 11112
rect 6880 11092 6882 11112
rect 6826 11056 6882 11092
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 2318 8744 2374 8800
rect 3422 8780 3424 8800
rect 3424 8780 3476 8800
rect 3476 8780 3478 8800
rect 3422 8744 3478 8780
rect 2134 7656 2190 7712
rect 2502 7404 2558 7440
rect 2502 7384 2504 7404
rect 2504 7384 2556 7404
rect 2556 7384 2558 7404
rect 3238 7404 3294 7440
rect 3238 7384 3240 7404
rect 3240 7384 3292 7404
rect 3292 7384 3294 7404
rect 938 4392 994 4448
rect 1306 3576 1362 3632
rect 2778 6024 2834 6080
rect 1858 5208 1914 5264
rect 1306 2760 1362 2816
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3974 6840 4030 6896
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3514 1944 3570 2000
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 1030 1164 1032 1184
rect 1032 1164 1084 1184
rect 1084 1164 1086 1184
rect 1030 1128 1086 1164
rect 6918 10668 6974 10704
rect 6918 10648 6920 10668
rect 6920 10648 6972 10668
rect 6972 10648 6974 10668
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 7654 11056 7710 11112
rect 8850 11192 8906 11248
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 7930 10376 7986 10432
rect 9218 11464 9274 11520
rect 8114 10240 8170 10296
rect 6918 8900 6974 8936
rect 6918 8880 6920 8900
rect 6920 8880 6972 8900
rect 6972 8880 6974 8900
rect 8022 10004 8024 10024
rect 8024 10004 8076 10024
rect 8076 10004 8078 10024
rect 8022 9968 8078 10004
rect 7838 8744 7894 8800
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8758 9868 8760 9888
rect 8760 9868 8812 9888
rect 8812 9868 8814 9888
rect 8758 9832 8814 9868
rect 9218 10376 9274 10432
rect 9034 10240 9090 10296
rect 9678 11736 9734 11792
rect 9678 11192 9734 11248
rect 9218 9596 9220 9616
rect 9220 9596 9272 9616
rect 9272 9596 9274 9616
rect 9218 9560 9274 9596
rect 9034 9424 9090 9480
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 9586 9868 9588 9888
rect 9588 9868 9640 9888
rect 9640 9868 9642 9888
rect 9586 9832 9642 9868
rect 9586 9580 9642 9616
rect 9586 9560 9588 9580
rect 9588 9560 9640 9580
rect 9640 9560 9642 9580
rect 10138 13368 10194 13424
rect 10138 12008 10194 12064
rect 10414 12008 10470 12064
rect 10046 11328 10102 11384
rect 9770 10376 9826 10432
rect 10414 11192 10470 11248
rect 10322 10512 10378 10568
rect 10138 10376 10194 10432
rect 10046 9968 10102 10024
rect 10322 9696 10378 9752
rect 10874 11192 10930 11248
rect 10966 10920 11022 10976
rect 11242 11328 11298 11384
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 11426 10648 11482 10704
rect 10782 10376 10838 10432
rect 9954 9560 10010 9616
rect 9678 8608 9734 8664
rect 9586 8492 9642 8528
rect 11150 10240 11206 10296
rect 10874 9424 10930 9480
rect 9954 8744 10010 8800
rect 9586 8472 9588 8492
rect 9588 8472 9640 8492
rect 9640 8472 9642 8492
rect 8758 8336 8814 8392
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 10138 8472 10194 8528
rect 10322 8472 10378 8528
rect 10782 8744 10838 8800
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 11794 11092 11796 11112
rect 11796 11092 11848 11112
rect 11848 11092 11850 11112
rect 11794 11056 11850 11092
rect 11978 11192 12034 11248
rect 11886 10648 11942 10704
rect 11886 10376 11942 10432
rect 12530 11600 12586 11656
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 12990 11756 13046 11792
rect 12990 11736 12992 11756
rect 12992 11736 13044 11756
rect 13044 11736 13046 11756
rect 12806 11600 12862 11656
rect 11886 9832 11942 9888
rect 11978 9696 12034 9752
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 13358 11192 13414 11248
rect 11610 9560 11666 9616
rect 11610 8336 11666 8392
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12530 9036 12586 9072
rect 12530 9016 12532 9036
rect 12532 9016 12584 9036
rect 12584 9016 12586 9036
rect 12070 8744 12126 8800
rect 12622 8744 12678 8800
rect 11242 7792 11298 7848
rect 11978 8336 12034 8392
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 13266 9424 13322 9480
rect 14002 11872 14058 11928
rect 13542 10920 13598 10976
rect 14186 10104 14242 10160
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 14186 9016 14242 9072
rect 15014 9832 15070 9888
rect 15382 10376 15438 10432
rect 14554 8744 14610 8800
rect 14462 8492 14518 8528
rect 14462 8472 14464 8492
rect 14464 8472 14516 8492
rect 14516 8472 14518 8492
rect 15198 8336 15254 8392
rect 15566 10104 15622 10160
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 15566 8472 15622 8528
rect 15566 8336 15622 8392
rect 16220 13082 16276 13084
rect 16300 13082 16356 13084
rect 16380 13082 16436 13084
rect 16460 13082 16516 13084
rect 16220 13030 16266 13082
rect 16266 13030 16276 13082
rect 16300 13030 16330 13082
rect 16330 13030 16342 13082
rect 16342 13030 16356 13082
rect 16380 13030 16394 13082
rect 16394 13030 16406 13082
rect 16406 13030 16436 13082
rect 16460 13030 16470 13082
rect 16470 13030 16516 13082
rect 16220 13028 16276 13030
rect 16300 13028 16356 13030
rect 16380 13028 16436 13030
rect 16460 13028 16516 13030
rect 16220 11994 16276 11996
rect 16300 11994 16356 11996
rect 16380 11994 16436 11996
rect 16460 11994 16516 11996
rect 16220 11942 16266 11994
rect 16266 11942 16276 11994
rect 16300 11942 16330 11994
rect 16330 11942 16342 11994
rect 16342 11942 16356 11994
rect 16380 11942 16394 11994
rect 16394 11942 16406 11994
rect 16406 11942 16436 11994
rect 16460 11942 16470 11994
rect 16470 11942 16516 11994
rect 16220 11940 16276 11942
rect 16300 11940 16356 11942
rect 16380 11940 16436 11942
rect 16460 11940 16516 11942
rect 16302 11092 16304 11112
rect 16304 11092 16356 11112
rect 16356 11092 16358 11112
rect 16302 11056 16358 11092
rect 16220 10906 16276 10908
rect 16300 10906 16356 10908
rect 16380 10906 16436 10908
rect 16460 10906 16516 10908
rect 16220 10854 16266 10906
rect 16266 10854 16276 10906
rect 16300 10854 16330 10906
rect 16330 10854 16342 10906
rect 16342 10854 16356 10906
rect 16380 10854 16394 10906
rect 16394 10854 16406 10906
rect 16406 10854 16436 10906
rect 16460 10854 16470 10906
rect 16470 10854 16516 10906
rect 16220 10852 16276 10854
rect 16300 10852 16356 10854
rect 16380 10852 16436 10854
rect 16460 10852 16516 10854
rect 16854 10648 16910 10704
rect 16220 9818 16276 9820
rect 16300 9818 16356 9820
rect 16380 9818 16436 9820
rect 16460 9818 16516 9820
rect 16220 9766 16266 9818
rect 16266 9766 16276 9818
rect 16300 9766 16330 9818
rect 16330 9766 16342 9818
rect 16342 9766 16356 9818
rect 16380 9766 16394 9818
rect 16394 9766 16406 9818
rect 16406 9766 16436 9818
rect 16460 9766 16470 9818
rect 16470 9766 16516 9818
rect 16220 9764 16276 9766
rect 16300 9764 16356 9766
rect 16380 9764 16436 9766
rect 16460 9764 16516 9766
rect 16220 8730 16276 8732
rect 16300 8730 16356 8732
rect 16380 8730 16436 8732
rect 16460 8730 16516 8732
rect 16220 8678 16266 8730
rect 16266 8678 16276 8730
rect 16300 8678 16330 8730
rect 16330 8678 16342 8730
rect 16342 8678 16356 8730
rect 16380 8678 16394 8730
rect 16394 8678 16406 8730
rect 16406 8678 16436 8730
rect 16460 8678 16470 8730
rect 16470 8678 16516 8730
rect 16220 8676 16276 8678
rect 16300 8676 16356 8678
rect 16380 8676 16436 8678
rect 16460 8676 16516 8678
rect 16210 7812 16266 7848
rect 16210 7792 16212 7812
rect 16212 7792 16264 7812
rect 16264 7792 16266 7812
rect 16220 7642 16276 7644
rect 16300 7642 16356 7644
rect 16380 7642 16436 7644
rect 16460 7642 16516 7644
rect 16220 7590 16266 7642
rect 16266 7590 16276 7642
rect 16300 7590 16330 7642
rect 16330 7590 16342 7642
rect 16342 7590 16356 7642
rect 16380 7590 16394 7642
rect 16394 7590 16406 7642
rect 16406 7590 16436 7642
rect 16460 7590 16470 7642
rect 16470 7590 16516 7642
rect 16220 7588 16276 7590
rect 16300 7588 16356 7590
rect 16380 7588 16436 7590
rect 16460 7588 16516 7590
rect 16220 6554 16276 6556
rect 16300 6554 16356 6556
rect 16380 6554 16436 6556
rect 16460 6554 16516 6556
rect 16220 6502 16266 6554
rect 16266 6502 16276 6554
rect 16300 6502 16330 6554
rect 16330 6502 16342 6554
rect 16342 6502 16356 6554
rect 16380 6502 16394 6554
rect 16394 6502 16406 6554
rect 16406 6502 16436 6554
rect 16460 6502 16470 6554
rect 16470 6502 16516 6554
rect 16220 6500 16276 6502
rect 16300 6500 16356 6502
rect 16380 6500 16436 6502
rect 16460 6500 16516 6502
rect 15842 6024 15898 6080
rect 16220 5466 16276 5468
rect 16300 5466 16356 5468
rect 16380 5466 16436 5468
rect 16460 5466 16516 5468
rect 16220 5414 16266 5466
rect 16266 5414 16276 5466
rect 16300 5414 16330 5466
rect 16330 5414 16342 5466
rect 16342 5414 16356 5466
rect 16380 5414 16394 5466
rect 16394 5414 16406 5466
rect 16406 5414 16436 5466
rect 16460 5414 16470 5466
rect 16470 5414 16516 5466
rect 16220 5412 16276 5414
rect 16300 5412 16356 5414
rect 16380 5412 16436 5414
rect 16460 5412 16516 5414
rect 17130 8916 17132 8936
rect 17132 8916 17184 8936
rect 17184 8916 17186 8936
rect 17130 8880 17186 8916
rect 16220 4378 16276 4380
rect 16300 4378 16356 4380
rect 16380 4378 16436 4380
rect 16460 4378 16516 4380
rect 16220 4326 16266 4378
rect 16266 4326 16276 4378
rect 16300 4326 16330 4378
rect 16330 4326 16342 4378
rect 16342 4326 16356 4378
rect 16380 4326 16394 4378
rect 16394 4326 16406 4378
rect 16406 4326 16436 4378
rect 16460 4326 16470 4378
rect 16470 4326 16516 4378
rect 16220 4324 16276 4326
rect 16300 4324 16356 4326
rect 16380 4324 16436 4326
rect 16460 4324 16516 4326
rect 15934 3576 15990 3632
rect 16220 3290 16276 3292
rect 16300 3290 16356 3292
rect 16380 3290 16436 3292
rect 16460 3290 16516 3292
rect 16220 3238 16266 3290
rect 16266 3238 16276 3290
rect 16300 3238 16330 3290
rect 16330 3238 16342 3290
rect 16342 3238 16356 3290
rect 16380 3238 16394 3290
rect 16394 3238 16406 3290
rect 16406 3238 16436 3290
rect 16460 3238 16470 3290
rect 16470 3238 16516 3290
rect 16220 3236 16276 3238
rect 16300 3236 16356 3238
rect 16380 3236 16436 3238
rect 16460 3236 16516 3238
rect 16220 2202 16276 2204
rect 16300 2202 16356 2204
rect 16380 2202 16436 2204
rect 16460 2202 16516 2204
rect 16220 2150 16266 2202
rect 16266 2150 16276 2202
rect 16300 2150 16330 2202
rect 16330 2150 16342 2202
rect 16342 2150 16356 2202
rect 16380 2150 16394 2202
rect 16394 2150 16406 2202
rect 16406 2150 16436 2202
rect 16460 2150 16470 2202
rect 16470 2150 16516 2202
rect 16220 2148 16276 2150
rect 16300 2148 16356 2150
rect 16380 2148 16436 2150
rect 16460 2148 16516 2150
rect 15382 1264 15438 1320
rect 16220 1114 16276 1116
rect 16300 1114 16356 1116
rect 16380 1114 16436 1116
rect 16460 1114 16516 1116
rect 16220 1062 16266 1114
rect 16266 1062 16276 1114
rect 16300 1062 16330 1114
rect 16330 1062 16342 1114
rect 16342 1062 16356 1114
rect 16380 1062 16394 1114
rect 16394 1062 16406 1114
rect 16406 1062 16436 1114
rect 16460 1062 16470 1114
rect 16470 1062 16516 1114
rect 16220 1060 16276 1062
rect 16300 1060 16356 1062
rect 16380 1060 16436 1062
rect 16460 1060 16516 1062
<< metal3 >>
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 12210 13632 12526 13633
rect 12210 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12526 13632
rect 12210 13567 12526 13568
rect 0 13426 800 13456
rect 3509 13426 3575 13429
rect 0 13424 3575 13426
rect 0 13368 3514 13424
rect 3570 13368 3575 13424
rect 0 13366 3575 13368
rect 0 13336 800 13366
rect 3509 13363 3575 13366
rect 10133 13426 10199 13429
rect 19200 13426 20000 13456
rect 10133 13424 20000 13426
rect 10133 13368 10138 13424
rect 10194 13368 20000 13424
rect 10133 13366 20000 13368
rect 10133 13363 10199 13366
rect 19200 13336 20000 13366
rect 8210 13088 8526 13089
rect 8210 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8526 13088
rect 8210 13023 8526 13024
rect 16210 13088 16526 13089
rect 16210 13024 16216 13088
rect 16280 13024 16296 13088
rect 16360 13024 16376 13088
rect 16440 13024 16456 13088
rect 16520 13024 16526 13088
rect 16210 13023 16526 13024
rect 0 12610 800 12640
rect 2129 12610 2195 12613
rect 0 12608 2195 12610
rect 0 12552 2134 12608
rect 2190 12552 2195 12608
rect 0 12550 2195 12552
rect 0 12520 800 12550
rect 2129 12547 2195 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12210 12544 12526 12545
rect 12210 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12526 12544
rect 12210 12479 12526 12480
rect 10133 12066 10199 12069
rect 10409 12066 10475 12069
rect 10133 12064 10475 12066
rect 10133 12008 10138 12064
rect 10194 12008 10414 12064
rect 10470 12008 10475 12064
rect 10133 12006 10475 12008
rect 10133 12003 10199 12006
rect 10409 12003 10475 12006
rect 8210 12000 8526 12001
rect 8210 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8526 12000
rect 8210 11935 8526 11936
rect 16210 12000 16526 12001
rect 16210 11936 16216 12000
rect 16280 11936 16296 12000
rect 16360 11936 16376 12000
rect 16440 11936 16456 12000
rect 16520 11936 16526 12000
rect 16210 11935 16526 11936
rect 9990 11868 9996 11932
rect 10060 11930 10066 11932
rect 13997 11930 14063 11933
rect 10060 11928 14063 11930
rect 10060 11872 14002 11928
rect 14058 11872 14063 11928
rect 10060 11870 14063 11872
rect 10060 11868 10066 11870
rect 13997 11867 14063 11870
rect 0 11794 800 11824
rect 3693 11794 3759 11797
rect 0 11792 3759 11794
rect 0 11736 3698 11792
rect 3754 11736 3759 11792
rect 0 11734 3759 11736
rect 0 11704 800 11734
rect 3693 11731 3759 11734
rect 9673 11794 9739 11797
rect 9806 11794 9812 11796
rect 9673 11792 9812 11794
rect 9673 11736 9678 11792
rect 9734 11736 9812 11792
rect 9673 11734 9812 11736
rect 9673 11731 9739 11734
rect 9806 11732 9812 11734
rect 9876 11732 9882 11796
rect 12985 11794 13051 11797
rect 11286 11792 13051 11794
rect 11286 11736 12990 11792
rect 13046 11736 13051 11792
rect 11286 11734 13051 11736
rect 9213 11522 9279 11525
rect 11286 11522 11346 11734
rect 12985 11731 13051 11734
rect 12525 11658 12591 11661
rect 12801 11658 12867 11661
rect 12525 11656 12867 11658
rect 12525 11600 12530 11656
rect 12586 11600 12806 11656
rect 12862 11600 12867 11656
rect 12525 11598 12867 11600
rect 12525 11595 12591 11598
rect 12801 11595 12867 11598
rect 9213 11520 11346 11522
rect 9213 11464 9218 11520
rect 9274 11464 11346 11520
rect 9213 11462 11346 11464
rect 9213 11459 9279 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 12210 11456 12526 11457
rect 12210 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12526 11456
rect 12210 11391 12526 11392
rect 10041 11386 10107 11389
rect 11237 11386 11303 11389
rect 10041 11384 11303 11386
rect 10041 11328 10046 11384
rect 10102 11328 11242 11384
rect 11298 11328 11303 11384
rect 10041 11326 11303 11328
rect 10041 11323 10107 11326
rect 11237 11323 11303 11326
rect 8845 11250 8911 11253
rect 4294 11248 8911 11250
rect 4294 11192 8850 11248
rect 8906 11192 8911 11248
rect 4294 11190 8911 11192
rect 0 10978 800 11008
rect 4294 10978 4354 11190
rect 8845 11187 8911 11190
rect 9673 11250 9739 11253
rect 9806 11250 9812 11252
rect 9673 11248 9812 11250
rect 9673 11192 9678 11248
rect 9734 11192 9812 11248
rect 9673 11190 9812 11192
rect 9673 11187 9739 11190
rect 9806 11188 9812 11190
rect 9876 11188 9882 11252
rect 10409 11250 10475 11253
rect 10869 11250 10935 11253
rect 10409 11248 10935 11250
rect 10409 11192 10414 11248
rect 10470 11192 10874 11248
rect 10930 11192 10935 11248
rect 10409 11190 10935 11192
rect 10409 11187 10475 11190
rect 10869 11187 10935 11190
rect 11973 11250 12039 11253
rect 13353 11250 13419 11253
rect 11973 11248 13419 11250
rect 11973 11192 11978 11248
rect 12034 11192 13358 11248
rect 13414 11192 13419 11248
rect 11973 11190 13419 11192
rect 11973 11187 12039 11190
rect 13353 11187 13419 11190
rect 6821 11114 6887 11117
rect 7649 11114 7715 11117
rect 11789 11114 11855 11117
rect 6821 11112 11855 11114
rect 6821 11056 6826 11112
rect 6882 11056 7654 11112
rect 7710 11056 11794 11112
rect 11850 11056 11855 11112
rect 6821 11054 11855 11056
rect 6821 11051 6887 11054
rect 7649 11051 7715 11054
rect 11789 11051 11855 11054
rect 16297 11114 16363 11117
rect 16297 11112 16682 11114
rect 16297 11056 16302 11112
rect 16358 11056 16682 11112
rect 16297 11054 16682 11056
rect 16297 11051 16363 11054
rect 0 10918 4354 10978
rect 10961 10978 11027 10981
rect 13537 10978 13603 10981
rect 10961 10976 13603 10978
rect 10961 10920 10966 10976
rect 11022 10920 13542 10976
rect 13598 10920 13603 10976
rect 10961 10918 13603 10920
rect 16622 10978 16682 11054
rect 19200 10978 20000 11008
rect 16622 10918 20000 10978
rect 0 10888 800 10918
rect 10961 10915 11027 10918
rect 13537 10915 13603 10918
rect 8210 10912 8526 10913
rect 8210 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8526 10912
rect 8210 10847 8526 10848
rect 16210 10912 16526 10913
rect 16210 10848 16216 10912
rect 16280 10848 16296 10912
rect 16360 10848 16376 10912
rect 16440 10848 16456 10912
rect 16520 10848 16526 10912
rect 19200 10888 20000 10918
rect 16210 10847 16526 10848
rect 2589 10706 2655 10709
rect 6913 10706 6979 10709
rect 11421 10706 11487 10709
rect 2589 10704 2790 10706
rect 2589 10648 2594 10704
rect 2650 10648 2790 10704
rect 2589 10646 2790 10648
rect 2589 10643 2655 10646
rect 2730 10570 2790 10646
rect 6913 10704 11487 10706
rect 6913 10648 6918 10704
rect 6974 10648 11426 10704
rect 11482 10648 11487 10704
rect 6913 10646 11487 10648
rect 6913 10643 6979 10646
rect 11421 10643 11487 10646
rect 11881 10706 11947 10709
rect 16849 10706 16915 10709
rect 11881 10704 16915 10706
rect 11881 10648 11886 10704
rect 11942 10648 16854 10704
rect 16910 10648 16915 10704
rect 11881 10646 16915 10648
rect 11881 10643 11947 10646
rect 16849 10643 16915 10646
rect 10317 10570 10383 10573
rect 2730 10568 10383 10570
rect 2730 10512 10322 10568
rect 10378 10512 10383 10568
rect 2730 10510 10383 10512
rect 10317 10507 10383 10510
rect 7925 10434 7991 10437
rect 9213 10434 9279 10437
rect 7925 10432 9279 10434
rect 7925 10376 7930 10432
rect 7986 10376 9218 10432
rect 9274 10376 9279 10432
rect 7925 10374 9279 10376
rect 7925 10371 7991 10374
rect 9213 10371 9279 10374
rect 9765 10434 9831 10437
rect 9990 10434 9996 10436
rect 9765 10432 9996 10434
rect 9765 10376 9770 10432
rect 9826 10376 9996 10432
rect 9765 10374 9996 10376
rect 9765 10371 9831 10374
rect 9990 10372 9996 10374
rect 10060 10372 10066 10436
rect 10133 10434 10199 10437
rect 10777 10434 10843 10437
rect 11881 10434 11947 10437
rect 10133 10432 11947 10434
rect 10133 10376 10138 10432
rect 10194 10376 10782 10432
rect 10838 10376 11886 10432
rect 11942 10376 11947 10432
rect 10133 10374 11947 10376
rect 10133 10371 10199 10374
rect 10777 10371 10843 10374
rect 11881 10371 11947 10374
rect 15377 10434 15443 10437
rect 15377 10432 15578 10434
rect 15377 10376 15382 10432
rect 15438 10376 15578 10432
rect 15377 10374 15578 10376
rect 15377 10371 15443 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12210 10368 12526 10369
rect 12210 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12526 10368
rect 12210 10303 12526 10304
rect 8109 10298 8175 10301
rect 9029 10298 9095 10301
rect 11145 10298 11211 10301
rect 8109 10296 11211 10298
rect 8109 10240 8114 10296
rect 8170 10240 9034 10296
rect 9090 10240 11150 10296
rect 11206 10240 11211 10296
rect 8109 10238 11211 10240
rect 8109 10235 8175 10238
rect 9029 10235 9095 10238
rect 11145 10235 11211 10238
rect 0 10162 800 10192
rect 15518 10165 15578 10374
rect 14181 10162 14247 10165
rect 0 10160 14247 10162
rect 0 10104 14186 10160
rect 14242 10104 14247 10160
rect 0 10102 14247 10104
rect 15518 10160 15627 10165
rect 15518 10104 15566 10160
rect 15622 10104 15627 10160
rect 15518 10102 15627 10104
rect 0 10072 800 10102
rect 14181 10099 14247 10102
rect 15561 10099 15627 10102
rect 8017 10026 8083 10029
rect 10041 10026 10107 10029
rect 8017 10024 10107 10026
rect 8017 9968 8022 10024
rect 8078 9968 10046 10024
rect 10102 9968 10107 10024
rect 8017 9966 10107 9968
rect 8017 9963 8083 9966
rect 10041 9963 10107 9966
rect 8753 9890 8819 9893
rect 9581 9890 9647 9893
rect 8753 9888 9647 9890
rect 8753 9832 8758 9888
rect 8814 9832 9586 9888
rect 9642 9832 9647 9888
rect 8753 9830 9647 9832
rect 8753 9827 8819 9830
rect 9581 9827 9647 9830
rect 11881 9890 11947 9893
rect 15009 9890 15075 9893
rect 11881 9888 15075 9890
rect 11881 9832 11886 9888
rect 11942 9832 15014 9888
rect 15070 9832 15075 9888
rect 11881 9830 15075 9832
rect 11881 9827 11947 9830
rect 15009 9827 15075 9830
rect 8210 9824 8526 9825
rect 8210 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8526 9824
rect 8210 9759 8526 9760
rect 16210 9824 16526 9825
rect 16210 9760 16216 9824
rect 16280 9760 16296 9824
rect 16360 9760 16376 9824
rect 16440 9760 16456 9824
rect 16520 9760 16526 9824
rect 16210 9759 16526 9760
rect 10317 9754 10383 9757
rect 11973 9754 12039 9757
rect 10317 9752 12039 9754
rect 10317 9696 10322 9752
rect 10378 9696 11978 9752
rect 12034 9696 12039 9752
rect 10317 9694 12039 9696
rect 10317 9691 10383 9694
rect 11973 9691 12039 9694
rect 9213 9618 9279 9621
rect 9581 9618 9647 9621
rect 9949 9618 10015 9621
rect 11605 9618 11671 9621
rect 9213 9616 9647 9618
rect 9213 9560 9218 9616
rect 9274 9560 9586 9616
rect 9642 9560 9647 9616
rect 9213 9558 9647 9560
rect 9213 9555 9279 9558
rect 9581 9555 9647 9558
rect 9768 9616 11671 9618
rect 9768 9560 9954 9616
rect 10010 9560 11610 9616
rect 11666 9560 11671 9616
rect 9768 9558 11671 9560
rect 9029 9482 9095 9485
rect 9768 9482 9828 9558
rect 9949 9555 10015 9558
rect 11605 9555 11671 9558
rect 9029 9480 9828 9482
rect 9029 9424 9034 9480
rect 9090 9424 9828 9480
rect 9029 9422 9828 9424
rect 10869 9482 10935 9485
rect 13261 9482 13327 9485
rect 10869 9480 13327 9482
rect 10869 9424 10874 9480
rect 10930 9424 13266 9480
rect 13322 9424 13327 9480
rect 10869 9422 13327 9424
rect 9029 9419 9095 9422
rect 10869 9419 10935 9422
rect 13261 9419 13327 9422
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12210 9280 12526 9281
rect 12210 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12526 9280
rect 12210 9215 12526 9216
rect 12525 9074 12591 9077
rect 14181 9074 14247 9077
rect 12525 9072 14247 9074
rect 12525 9016 12530 9072
rect 12586 9016 14186 9072
rect 14242 9016 14247 9072
rect 12525 9014 14247 9016
rect 12525 9011 12591 9014
rect 14181 9011 14247 9014
rect 6913 8938 6979 8941
rect 17125 8938 17191 8941
rect 6913 8936 17191 8938
rect 6913 8880 6918 8936
rect 6974 8880 17130 8936
rect 17186 8880 17191 8936
rect 6913 8878 17191 8880
rect 6913 8875 6979 8878
rect 17125 8875 17191 8878
rect 2313 8802 2379 8805
rect 3417 8802 3483 8805
rect 7833 8802 7899 8805
rect 2313 8800 7899 8802
rect 2313 8744 2318 8800
rect 2374 8744 3422 8800
rect 3478 8744 7838 8800
rect 7894 8744 7899 8800
rect 2313 8742 7899 8744
rect 2313 8739 2379 8742
rect 3417 8739 3483 8742
rect 7833 8739 7899 8742
rect 9949 8802 10015 8805
rect 10777 8802 10843 8805
rect 9949 8800 10843 8802
rect 9949 8744 9954 8800
rect 10010 8744 10782 8800
rect 10838 8744 10843 8800
rect 9949 8742 10843 8744
rect 9949 8739 10015 8742
rect 10777 8739 10843 8742
rect 12065 8802 12131 8805
rect 12617 8802 12683 8805
rect 14549 8802 14615 8805
rect 12065 8800 14615 8802
rect 12065 8744 12070 8800
rect 12126 8744 12622 8800
rect 12678 8744 14554 8800
rect 14610 8744 14615 8800
rect 12065 8742 14615 8744
rect 12065 8739 12131 8742
rect 12617 8739 12683 8742
rect 14549 8739 14615 8742
rect 8210 8736 8526 8737
rect 8210 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8526 8736
rect 8210 8671 8526 8672
rect 16210 8736 16526 8737
rect 16210 8672 16216 8736
rect 16280 8672 16296 8736
rect 16360 8672 16376 8736
rect 16440 8672 16456 8736
rect 16520 8672 16526 8736
rect 16210 8671 16526 8672
rect 9673 8666 9739 8669
rect 9673 8664 10380 8666
rect 9673 8608 9678 8664
rect 9734 8608 10380 8664
rect 9673 8606 10380 8608
rect 9673 8603 9739 8606
rect 0 8530 800 8560
rect 10320 8533 10380 8606
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 800 8470
rect 1209 8467 1275 8470
rect 9581 8530 9647 8533
rect 10133 8530 10199 8533
rect 9581 8528 10199 8530
rect 9581 8472 9586 8528
rect 9642 8472 10138 8528
rect 10194 8472 10199 8528
rect 9581 8470 10199 8472
rect 9581 8467 9647 8470
rect 10133 8467 10199 8470
rect 10317 8528 10383 8533
rect 10317 8472 10322 8528
rect 10378 8472 10383 8528
rect 10317 8467 10383 8472
rect 14457 8530 14523 8533
rect 15561 8530 15627 8533
rect 19200 8530 20000 8560
rect 14457 8528 15394 8530
rect 14457 8472 14462 8528
rect 14518 8472 15394 8528
rect 14457 8470 15394 8472
rect 14457 8467 14523 8470
rect 8753 8394 8819 8397
rect 11605 8394 11671 8397
rect 8753 8392 11671 8394
rect 8753 8336 8758 8392
rect 8814 8336 11610 8392
rect 11666 8336 11671 8392
rect 8753 8334 11671 8336
rect 8753 8331 8819 8334
rect 11605 8331 11671 8334
rect 11973 8394 12039 8397
rect 15193 8394 15259 8397
rect 11973 8392 15259 8394
rect 11973 8336 11978 8392
rect 12034 8336 15198 8392
rect 15254 8336 15259 8392
rect 11973 8334 15259 8336
rect 15334 8394 15394 8470
rect 15561 8528 20000 8530
rect 15561 8472 15566 8528
rect 15622 8472 20000 8528
rect 15561 8470 20000 8472
rect 15561 8467 15627 8470
rect 19200 8440 20000 8470
rect 15561 8394 15627 8397
rect 15334 8392 15627 8394
rect 15334 8336 15566 8392
rect 15622 8336 15627 8392
rect 15334 8334 15627 8336
rect 11973 8331 12039 8334
rect 15193 8331 15259 8334
rect 15561 8331 15627 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 12210 8192 12526 8193
rect 12210 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12526 8192
rect 12210 8127 12526 8128
rect 11237 7850 11303 7853
rect 16205 7850 16271 7853
rect 11237 7848 16271 7850
rect 11237 7792 11242 7848
rect 11298 7792 16210 7848
rect 16266 7792 16271 7848
rect 11237 7790 16271 7792
rect 11237 7787 11303 7790
rect 16205 7787 16271 7790
rect 0 7714 800 7744
rect 2129 7714 2195 7717
rect 0 7712 2195 7714
rect 0 7656 2134 7712
rect 2190 7656 2195 7712
rect 0 7654 2195 7656
rect 0 7624 800 7654
rect 2129 7651 2195 7654
rect 8210 7648 8526 7649
rect 8210 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8526 7648
rect 8210 7583 8526 7584
rect 16210 7648 16526 7649
rect 16210 7584 16216 7648
rect 16280 7584 16296 7648
rect 16360 7584 16376 7648
rect 16440 7584 16456 7648
rect 16520 7584 16526 7648
rect 16210 7583 16526 7584
rect 2497 7442 2563 7445
rect 3233 7442 3299 7445
rect 2497 7440 3299 7442
rect 2497 7384 2502 7440
rect 2558 7384 3238 7440
rect 3294 7384 3299 7440
rect 2497 7382 3299 7384
rect 2497 7379 2563 7382
rect 3233 7379 3299 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12210 7104 12526 7105
rect 12210 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12526 7104
rect 12210 7039 12526 7040
rect 0 6898 800 6928
rect 3969 6898 4035 6901
rect 0 6896 4035 6898
rect 0 6840 3974 6896
rect 4030 6840 4035 6896
rect 0 6838 4035 6840
rect 0 6808 800 6838
rect 3969 6835 4035 6838
rect 8210 6560 8526 6561
rect 8210 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8526 6560
rect 8210 6495 8526 6496
rect 16210 6560 16526 6561
rect 16210 6496 16216 6560
rect 16280 6496 16296 6560
rect 16360 6496 16376 6560
rect 16440 6496 16456 6560
rect 16520 6496 16526 6560
rect 16210 6495 16526 6496
rect 0 6082 800 6112
rect 2773 6082 2839 6085
rect 0 6080 2839 6082
rect 0 6024 2778 6080
rect 2834 6024 2839 6080
rect 0 6022 2839 6024
rect 0 5992 800 6022
rect 2773 6019 2839 6022
rect 15837 6082 15903 6085
rect 19200 6082 20000 6112
rect 15837 6080 20000 6082
rect 15837 6024 15842 6080
rect 15898 6024 20000 6080
rect 15837 6022 20000 6024
rect 15837 6019 15903 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12210 6016 12526 6017
rect 12210 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12526 6016
rect 19200 5992 20000 6022
rect 12210 5951 12526 5952
rect 8210 5472 8526 5473
rect 8210 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8526 5472
rect 8210 5407 8526 5408
rect 16210 5472 16526 5473
rect 16210 5408 16216 5472
rect 16280 5408 16296 5472
rect 16360 5408 16376 5472
rect 16440 5408 16456 5472
rect 16520 5408 16526 5472
rect 16210 5407 16526 5408
rect 0 5266 800 5296
rect 1853 5266 1919 5269
rect 0 5264 1919 5266
rect 0 5208 1858 5264
rect 1914 5208 1919 5264
rect 0 5206 1919 5208
rect 0 5176 800 5206
rect 1853 5203 1919 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12210 4928 12526 4929
rect 12210 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12526 4928
rect 12210 4863 12526 4864
rect 0 4450 800 4480
rect 933 4450 999 4453
rect 0 4448 999 4450
rect 0 4392 938 4448
rect 994 4392 999 4448
rect 0 4390 999 4392
rect 0 4360 800 4390
rect 933 4387 999 4390
rect 8210 4384 8526 4385
rect 8210 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8526 4384
rect 8210 4319 8526 4320
rect 16210 4384 16526 4385
rect 16210 4320 16216 4384
rect 16280 4320 16296 4384
rect 16360 4320 16376 4384
rect 16440 4320 16456 4384
rect 16520 4320 16526 4384
rect 16210 4319 16526 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12210 3840 12526 3841
rect 12210 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12526 3840
rect 12210 3775 12526 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 15929 3634 15995 3637
rect 19200 3634 20000 3664
rect 15929 3632 20000 3634
rect 15929 3576 15934 3632
rect 15990 3576 20000 3632
rect 15929 3574 20000 3576
rect 15929 3571 15995 3574
rect 19200 3544 20000 3574
rect 8210 3296 8526 3297
rect 8210 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8526 3296
rect 8210 3231 8526 3232
rect 16210 3296 16526 3297
rect 16210 3232 16216 3296
rect 16280 3232 16296 3296
rect 16360 3232 16376 3296
rect 16440 3232 16456 3296
rect 16520 3232 16526 3296
rect 16210 3231 16526 3232
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12210 2752 12526 2753
rect 12210 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12526 2752
rect 12210 2687 12526 2688
rect 8210 2208 8526 2209
rect 8210 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8526 2208
rect 8210 2143 8526 2144
rect 16210 2208 16526 2209
rect 16210 2144 16216 2208
rect 16280 2144 16296 2208
rect 16360 2144 16376 2208
rect 16440 2144 16456 2208
rect 16520 2144 16526 2208
rect 16210 2143 16526 2144
rect 0 2002 800 2032
rect 3509 2002 3575 2005
rect 0 2000 3575 2002
rect 0 1944 3514 2000
rect 3570 1944 3575 2000
rect 0 1942 3575 1944
rect 0 1912 800 1942
rect 3509 1939 3575 1942
rect 4210 1664 4526 1665
rect 4210 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4526 1664
rect 4210 1599 4526 1600
rect 12210 1664 12526 1665
rect 12210 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12526 1664
rect 12210 1599 12526 1600
rect 15377 1322 15443 1325
rect 15377 1320 17970 1322
rect 15377 1264 15382 1320
rect 15438 1264 17970 1320
rect 15377 1262 17970 1264
rect 15377 1259 15443 1262
rect 0 1186 800 1216
rect 1025 1186 1091 1189
rect 0 1184 1091 1186
rect 0 1128 1030 1184
rect 1086 1128 1091 1184
rect 0 1126 1091 1128
rect 17910 1186 17970 1262
rect 19200 1186 20000 1216
rect 17910 1126 20000 1186
rect 0 1096 800 1126
rect 1025 1123 1091 1126
rect 8210 1120 8526 1121
rect 8210 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8526 1120
rect 8210 1055 8526 1056
rect 16210 1120 16526 1121
rect 16210 1056 16216 1120
rect 16280 1056 16296 1120
rect 16360 1056 16376 1120
rect 16440 1056 16456 1120
rect 16520 1056 16526 1120
rect 19200 1096 20000 1126
rect 16210 1055 16526 1056
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 16216 13084 16280 13088
rect 16216 13028 16220 13084
rect 16220 13028 16276 13084
rect 16276 13028 16280 13084
rect 16216 13024 16280 13028
rect 16296 13084 16360 13088
rect 16296 13028 16300 13084
rect 16300 13028 16356 13084
rect 16356 13028 16360 13084
rect 16296 13024 16360 13028
rect 16376 13084 16440 13088
rect 16376 13028 16380 13084
rect 16380 13028 16436 13084
rect 16436 13028 16440 13084
rect 16376 13024 16440 13028
rect 16456 13084 16520 13088
rect 16456 13028 16460 13084
rect 16460 13028 16516 13084
rect 16516 13028 16520 13084
rect 16456 13024 16520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 16216 11996 16280 12000
rect 16216 11940 16220 11996
rect 16220 11940 16276 11996
rect 16276 11940 16280 11996
rect 16216 11936 16280 11940
rect 16296 11996 16360 12000
rect 16296 11940 16300 11996
rect 16300 11940 16356 11996
rect 16356 11940 16360 11996
rect 16296 11936 16360 11940
rect 16376 11996 16440 12000
rect 16376 11940 16380 11996
rect 16380 11940 16436 11996
rect 16436 11940 16440 11996
rect 16376 11936 16440 11940
rect 16456 11996 16520 12000
rect 16456 11940 16460 11996
rect 16460 11940 16516 11996
rect 16516 11940 16520 11996
rect 16456 11936 16520 11940
rect 9996 11868 10060 11932
rect 9812 11732 9876 11796
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 9812 11188 9876 11252
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 16216 10908 16280 10912
rect 16216 10852 16220 10908
rect 16220 10852 16276 10908
rect 16276 10852 16280 10908
rect 16216 10848 16280 10852
rect 16296 10908 16360 10912
rect 16296 10852 16300 10908
rect 16300 10852 16356 10908
rect 16356 10852 16360 10908
rect 16296 10848 16360 10852
rect 16376 10908 16440 10912
rect 16376 10852 16380 10908
rect 16380 10852 16436 10908
rect 16436 10852 16440 10908
rect 16376 10848 16440 10852
rect 16456 10908 16520 10912
rect 16456 10852 16460 10908
rect 16460 10852 16516 10908
rect 16516 10852 16520 10908
rect 16456 10848 16520 10852
rect 9996 10372 10060 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 16216 9820 16280 9824
rect 16216 9764 16220 9820
rect 16220 9764 16276 9820
rect 16276 9764 16280 9820
rect 16216 9760 16280 9764
rect 16296 9820 16360 9824
rect 16296 9764 16300 9820
rect 16300 9764 16356 9820
rect 16356 9764 16360 9820
rect 16296 9760 16360 9764
rect 16376 9820 16440 9824
rect 16376 9764 16380 9820
rect 16380 9764 16436 9820
rect 16436 9764 16440 9820
rect 16376 9760 16440 9764
rect 16456 9820 16520 9824
rect 16456 9764 16460 9820
rect 16460 9764 16516 9820
rect 16516 9764 16520 9820
rect 16456 9760 16520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 16216 8732 16280 8736
rect 16216 8676 16220 8732
rect 16220 8676 16276 8732
rect 16276 8676 16280 8732
rect 16216 8672 16280 8676
rect 16296 8732 16360 8736
rect 16296 8676 16300 8732
rect 16300 8676 16356 8732
rect 16356 8676 16360 8732
rect 16296 8672 16360 8676
rect 16376 8732 16440 8736
rect 16376 8676 16380 8732
rect 16380 8676 16436 8732
rect 16436 8676 16440 8732
rect 16376 8672 16440 8676
rect 16456 8732 16520 8736
rect 16456 8676 16460 8732
rect 16460 8676 16516 8732
rect 16516 8676 16520 8732
rect 16456 8672 16520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 16216 7644 16280 7648
rect 16216 7588 16220 7644
rect 16220 7588 16276 7644
rect 16276 7588 16280 7644
rect 16216 7584 16280 7588
rect 16296 7644 16360 7648
rect 16296 7588 16300 7644
rect 16300 7588 16356 7644
rect 16356 7588 16360 7644
rect 16296 7584 16360 7588
rect 16376 7644 16440 7648
rect 16376 7588 16380 7644
rect 16380 7588 16436 7644
rect 16436 7588 16440 7644
rect 16376 7584 16440 7588
rect 16456 7644 16520 7648
rect 16456 7588 16460 7644
rect 16460 7588 16516 7644
rect 16516 7588 16520 7644
rect 16456 7584 16520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 16216 6556 16280 6560
rect 16216 6500 16220 6556
rect 16220 6500 16276 6556
rect 16276 6500 16280 6556
rect 16216 6496 16280 6500
rect 16296 6556 16360 6560
rect 16296 6500 16300 6556
rect 16300 6500 16356 6556
rect 16356 6500 16360 6556
rect 16296 6496 16360 6500
rect 16376 6556 16440 6560
rect 16376 6500 16380 6556
rect 16380 6500 16436 6556
rect 16436 6500 16440 6556
rect 16376 6496 16440 6500
rect 16456 6556 16520 6560
rect 16456 6500 16460 6556
rect 16460 6500 16516 6556
rect 16516 6500 16520 6556
rect 16456 6496 16520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 16216 5468 16280 5472
rect 16216 5412 16220 5468
rect 16220 5412 16276 5468
rect 16276 5412 16280 5468
rect 16216 5408 16280 5412
rect 16296 5468 16360 5472
rect 16296 5412 16300 5468
rect 16300 5412 16356 5468
rect 16356 5412 16360 5468
rect 16296 5408 16360 5412
rect 16376 5468 16440 5472
rect 16376 5412 16380 5468
rect 16380 5412 16436 5468
rect 16436 5412 16440 5468
rect 16376 5408 16440 5412
rect 16456 5468 16520 5472
rect 16456 5412 16460 5468
rect 16460 5412 16516 5468
rect 16516 5412 16520 5468
rect 16456 5408 16520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 16216 4380 16280 4384
rect 16216 4324 16220 4380
rect 16220 4324 16276 4380
rect 16276 4324 16280 4380
rect 16216 4320 16280 4324
rect 16296 4380 16360 4384
rect 16296 4324 16300 4380
rect 16300 4324 16356 4380
rect 16356 4324 16360 4380
rect 16296 4320 16360 4324
rect 16376 4380 16440 4384
rect 16376 4324 16380 4380
rect 16380 4324 16436 4380
rect 16436 4324 16440 4380
rect 16376 4320 16440 4324
rect 16456 4380 16520 4384
rect 16456 4324 16460 4380
rect 16460 4324 16516 4380
rect 16516 4324 16520 4380
rect 16456 4320 16520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 16216 3292 16280 3296
rect 16216 3236 16220 3292
rect 16220 3236 16276 3292
rect 16276 3236 16280 3292
rect 16216 3232 16280 3236
rect 16296 3292 16360 3296
rect 16296 3236 16300 3292
rect 16300 3236 16356 3292
rect 16356 3236 16360 3292
rect 16296 3232 16360 3236
rect 16376 3292 16440 3296
rect 16376 3236 16380 3292
rect 16380 3236 16436 3292
rect 16436 3236 16440 3292
rect 16376 3232 16440 3236
rect 16456 3292 16520 3296
rect 16456 3236 16460 3292
rect 16460 3236 16516 3292
rect 16516 3236 16520 3292
rect 16456 3232 16520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 16216 2204 16280 2208
rect 16216 2148 16220 2204
rect 16220 2148 16276 2204
rect 16276 2148 16280 2204
rect 16216 2144 16280 2148
rect 16296 2204 16360 2208
rect 16296 2148 16300 2204
rect 16300 2148 16356 2204
rect 16356 2148 16360 2204
rect 16296 2144 16360 2148
rect 16376 2204 16440 2208
rect 16376 2148 16380 2204
rect 16380 2148 16436 2204
rect 16436 2148 16440 2204
rect 16376 2144 16440 2148
rect 16456 2204 16520 2208
rect 16456 2148 16460 2204
rect 16460 2148 16516 2204
rect 16516 2148 16520 2204
rect 16456 2144 16520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
rect 16216 1116 16280 1120
rect 16216 1060 16220 1116
rect 16220 1060 16276 1116
rect 16276 1060 16280 1116
rect 16216 1056 16280 1060
rect 16296 1116 16360 1120
rect 16296 1060 16300 1116
rect 16300 1060 16356 1116
rect 16356 1060 16360 1116
rect 16296 1056 16360 1060
rect 16376 1116 16440 1120
rect 16376 1060 16380 1116
rect 16380 1060 16436 1116
rect 16436 1060 16440 1116
rect 16376 1056 16440 1060
rect 16456 1116 16520 1120
rect 16456 1060 16460 1116
rect 16460 1060 16516 1116
rect 16516 1060 16520 1116
rect 16456 1056 16520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12528 12544
rect 9995 11932 10061 11933
rect 9995 11868 9996 11932
rect 10060 11868 10061 11932
rect 9995 11867 10061 11868
rect 9811 11796 9877 11797
rect 9811 11732 9812 11796
rect 9876 11732 9877 11796
rect 9811 11731 9877 11732
rect 9814 11253 9874 11731
rect 9811 11252 9877 11253
rect 9811 11188 9812 11252
rect 9876 11188 9877 11252
rect 9811 11187 9877 11188
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 9998 10437 10058 11867
rect 12208 11456 12528 12480
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 9995 10436 10061 10437
rect 9995 10372 9996 10436
rect 10060 10372 10061 10436
rect 9995 10371 10061 10372
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 7648 8528 8672
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 3840 12528 4864
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
rect 16208 13088 16528 13648
rect 16208 13024 16216 13088
rect 16280 13024 16296 13088
rect 16360 13024 16376 13088
rect 16440 13024 16456 13088
rect 16520 13024 16528 13088
rect 16208 12000 16528 13024
rect 16208 11936 16216 12000
rect 16280 11936 16296 12000
rect 16360 11936 16376 12000
rect 16440 11936 16456 12000
rect 16520 11936 16528 12000
rect 16208 10912 16528 11936
rect 16208 10848 16216 10912
rect 16280 10848 16296 10912
rect 16360 10848 16376 10912
rect 16440 10848 16456 10912
rect 16520 10848 16528 10912
rect 16208 9824 16528 10848
rect 16208 9760 16216 9824
rect 16280 9760 16296 9824
rect 16360 9760 16376 9824
rect 16440 9760 16456 9824
rect 16520 9760 16528 9824
rect 16208 8736 16528 9760
rect 16208 8672 16216 8736
rect 16280 8672 16296 8736
rect 16360 8672 16376 8736
rect 16440 8672 16456 8736
rect 16520 8672 16528 8736
rect 16208 7648 16528 8672
rect 16208 7584 16216 7648
rect 16280 7584 16296 7648
rect 16360 7584 16376 7648
rect 16440 7584 16456 7648
rect 16520 7584 16528 7648
rect 16208 6560 16528 7584
rect 16208 6496 16216 6560
rect 16280 6496 16296 6560
rect 16360 6496 16376 6560
rect 16440 6496 16456 6560
rect 16520 6496 16528 6560
rect 16208 5472 16528 6496
rect 16208 5408 16216 5472
rect 16280 5408 16296 5472
rect 16360 5408 16376 5472
rect 16440 5408 16456 5472
rect 16520 5408 16528 5472
rect 16208 4384 16528 5408
rect 16208 4320 16216 4384
rect 16280 4320 16296 4384
rect 16360 4320 16376 4384
rect 16440 4320 16456 4384
rect 16520 4320 16528 4384
rect 16208 3296 16528 4320
rect 16208 3232 16216 3296
rect 16280 3232 16296 3296
rect 16360 3232 16376 3296
rect 16440 3232 16456 3296
rect 16520 3232 16528 3296
rect 16208 2208 16528 3232
rect 16208 2144 16216 2208
rect 16280 2144 16296 2208
rect 16360 2144 16376 2208
rect 16440 2144 16456 2208
rect 16520 2144 16528 2208
rect 16208 1120 16528 2144
rect 16208 1056 16216 1120
rect 16280 1056 16296 1120
rect 16360 1056 16376 1120
rect 16440 1056 16456 1120
rect 16520 1056 16528 1120
rect 16208 1040 16528 1056
use sky130_fd_sc_hd__inv_2  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1683767628
transform 1 0 9016 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1683767628
transform 1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1683767628
transform 1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1683767628
transform 1 0 11592 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1683767628
transform 1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1683767628
transform 1 0 1564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1683767628
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 15456 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2760 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _192_
timestamp 1683767628
transform 1 0 6440 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1683767628
transform 1 0 10488 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _194_
timestamp 1683767628
transform 1 0 4876 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1683767628
transform 1 0 2576 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3956 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1683767628
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 6532 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _201_
timestamp 1683767628
transform 1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _202_
timestamp 1683767628
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 6808 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _204_
timestamp 1683767628
transform 1 0 6624 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _205_
timestamp 1683767628
transform 1 0 5428 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _206_
timestamp 1683767628
transform 1 0 3036 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 1683767628
transform 1 0 3864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4692 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5428 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4600 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _212_
timestamp 1683767628
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _213_
timestamp 1683767628
transform 1 0 4784 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2116 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _215_
timestamp 1683767628
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _216_
timestamp 1683767628
transform 1 0 5152 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _217_
timestamp 1683767628
transform 1 0 5428 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3956 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _219_
timestamp 1683767628
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _220_
timestamp 1683767628
transform 1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2392 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _222_
timestamp 1683767628
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _223_
timestamp 1683767628
transform 1 0 2944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _224_
timestamp 1683767628
transform 1 0 4600 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _225_
timestamp 1683767628
transform 1 0 1656 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _226_
timestamp 1683767628
transform 1 0 1748 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _227_
timestamp 1683767628
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1683767628
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1840 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _232_
timestamp 1683767628
transform 1 0 3036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2024 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 1683767628
transform 1 0 10580 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _236_
timestamp 1683767628
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _237_
timestamp 1683767628
transform 1 0 12420 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1683767628
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _239_
timestamp 1683767628
transform 1 0 12880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _240_
timestamp 1683767628
transform 1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _241_
timestamp 1683767628
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _242_
timestamp 1683767628
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1683767628
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _244_
timestamp 1683767628
transform 1 0 6624 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 16376 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _247_
timestamp 1683767628
transform 1 0 2116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_1  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2300 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 7544 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _250_
timestamp 1683767628
transform 1 0 9568 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _251_
timestamp 1683767628
transform 1 0 8648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _252_
timestamp 1683767628
transform 1 0 11408 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 7268 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _254_
timestamp 1683767628
transform 1 0 7452 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp 1683767628
transform 1 0 11684 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _256_
timestamp 1683767628
transform 1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _257_
timestamp 1683767628
transform 1 0 12972 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _258_
timestamp 1683767628
transform 1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _259_
timestamp 1683767628
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _260_
timestamp 1683767628
transform 1 0 8372 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _261_
timestamp 1683767628
transform 1 0 10304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 9384 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _263_
timestamp 1683767628
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _264_
timestamp 1683767628
transform 1 0 11316 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _265_
timestamp 1683767628
transform 1 0 12512 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _266_
timestamp 1683767628
transform 1 0 12696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12512 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _268_
timestamp 1683767628
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _269_
timestamp 1683767628
transform 1 0 13708 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1683767628
transform 1 0 14168 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _271_
timestamp 1683767628
transform 1 0 14168 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _272_
timestamp 1683767628
transform 1 0 14076 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1683767628
transform 1 0 10304 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _274_
timestamp 1683767628
transform 1 0 11592 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _275_
timestamp 1683767628
transform 1 0 10120 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _276_
timestamp 1683767628
transform 1 0 10028 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 9292 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _278_
timestamp 1683767628
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _279_
timestamp 1683767628
transform 1 0 6164 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1683767628
transform 1 0 7360 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1683767628
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8648 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _283_
timestamp 1683767628
transform 1 0 8464 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _284_
timestamp 1683767628
transform 1 0 9476 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _285_
timestamp 1683767628
transform 1 0 7636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _286_
timestamp 1683767628
transform 1 0 9476 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _287_
timestamp 1683767628
transform 1 0 9200 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 1683767628
transform 1 0 10672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _289_
timestamp 1683767628
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _290_
timestamp 1683767628
transform 1 0 9016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _291_
timestamp 1683767628
transform 1 0 10120 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _292_
timestamp 1683767628
transform 1 0 7452 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 9292 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 6440 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1683767628
transform 1 0 16744 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _296_
timestamp 1683767628
transform 1 0 17296 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _297_
timestamp 1683767628
transform 1 0 16928 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _298_
timestamp 1683767628
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _299_
timestamp 1683767628
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp 1683767628
transform 1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 7452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1683767628
transform 1 0 13064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _303_
timestamp 1683767628
transform 1 0 14260 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _304_
timestamp 1683767628
transform 1 0 10672 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8280 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1683767628
transform 1 0 9016 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10120 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 11500 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _309_
timestamp 1683767628
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _310_
timestamp 1683767628
transform 1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _311_
timestamp 1683767628
transform 1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _312_
timestamp 1683767628
transform 1 0 14352 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _313_
timestamp 1683767628
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _314_
timestamp 1683767628
transform 1 0 9936 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _315_
timestamp 1683767628
transform 1 0 8464 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _316_
timestamp 1683767628
transform 1 0 10580 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _317_
timestamp 1683767628
transform 1 0 4232 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _318_
timestamp 1683767628
transform 1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _319_
timestamp 1683767628
transform 1 0 9568 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _320_
timestamp 1683767628
transform 1 0 1656 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _321_
timestamp 1683767628
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _322_
timestamp 1683767628
transform 1 0 7544 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _323_
timestamp 1683767628
transform 1 0 6624 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _324_
timestamp 1683767628
transform 1 0 6532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10488 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _326_
timestamp 1683767628
transform 1 0 10396 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _327_
timestamp 1683767628
transform 1 0 10488 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _328_
timestamp 1683767628
transform 1 0 5520 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _329_
timestamp 1683767628
transform 1 0 6900 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 1683767628
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _331_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 7912 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _332_
timestamp 1683767628
transform 1 0 7636 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _333_
timestamp 1683767628
transform 1 0 7360 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _334_
timestamp 1683767628
transform 1 0 6164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _335_
timestamp 1683767628
transform 1 0 8832 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _336_
timestamp 1683767628
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _337_
timestamp 1683767628
transform 1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _338_
timestamp 1683767628
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _339_
timestamp 1683767628
transform 1 0 6900 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _340_
timestamp 1683767628
transform 1 0 6532 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _341_
timestamp 1683767628
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _342_
timestamp 1683767628
transform 1 0 12236 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _343_
timestamp 1683767628
transform 1 0 9016 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _344_
timestamp 1683767628
transform 1 0 8648 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _345_
timestamp 1683767628
transform 1 0 9476 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _346_
timestamp 1683767628
transform 1 0 11776 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _347_
timestamp 1683767628
transform 1 0 12236 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _348_
timestamp 1683767628
transform 1 0 13064 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _349_
timestamp 1683767628
transform 1 0 13064 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _350_
timestamp 1683767628
transform 1 0 15548 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _351_
timestamp 1683767628
transform 1 0 13340 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _352_
timestamp 1683767628
transform 1 0 15824 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _353_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _354_
timestamp 1683767628
transform 1 0 14536 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _355_
timestamp 1683767628
transform 1 0 11868 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _356_
timestamp 1683767628
transform 1 0 12604 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _357_
timestamp 1683767628
transform 1 0 9752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _358_
timestamp 1683767628
transform 1 0 10120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _359_
timestamp 1683767628
transform 1 0 9476 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _360_
timestamp 1683767628
transform 1 0 12420 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _361_
timestamp 1683767628
transform 1 0 15548 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _362_
timestamp 1683767628
transform 1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _363_
timestamp 1683767628
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _364_
timestamp 1683767628
transform 1 0 15824 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _365_
timestamp 1683767628
transform 1 0 15732 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _366_
timestamp 1683767628
transform 1 0 14904 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _367_
timestamp 1683767628
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _368_
timestamp 1683767628
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _369_
timestamp 1683767628
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _370_
timestamp 1683767628
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _371_
timestamp 1683767628
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _372_
timestamp 1683767628
transform 1 0 10948 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _373_
timestamp 1683767628
transform 1 0 10764 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _374_
timestamp 1683767628
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1683767628
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _376_
timestamp 1683767628
transform 1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _377_
timestamp 1683767628
transform 1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _378_
timestamp 1683767628
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _379_
timestamp 1683767628
transform 1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _380_
timestamp 1683767628
transform 1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _381_
timestamp 1683767628
transform 1 0 16744 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _382_
timestamp 1683767628
transform 1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _383_
timestamp 1683767628
transform 1 0 11868 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _384_
timestamp 1683767628
transform 1 0 14168 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _385_
timestamp 1683767628
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _386_
timestamp 1683767628
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _387_
timestamp 1683767628
transform 1 0 4232 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _388_
timestamp 1683767628
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _389_
timestamp 1683767628
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _390_
timestamp 1683767628
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 13892 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _392_
timestamp 1683767628
transform 1 0 14168 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _393_
timestamp 1683767628
transform 1 0 13800 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _394_
timestamp 1683767628
transform 1 0 6440 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _395_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8372 0 -1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1683767628
transform 1 0 9844 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10120 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _398_
timestamp 1683767628
transform 1 0 7176 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1683767628
transform 1 0 9016 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1683767628
transform 1 0 6808 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _401_
timestamp 1683767628
transform 1 0 9292 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1683767628
transform 1 0 11592 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1683767628
transform 1 0 14168 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _404_
timestamp 1683767628
transform 1 0 14168 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _405_
timestamp 1683767628
transform 1 0 13708 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _406_
timestamp 1683767628
transform 1 0 11684 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _407_
timestamp 1683767628
transform 1 0 13708 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _408_
timestamp 1683767628
transform 1 0 14168 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _409_
timestamp 1683767628
transform 1 0 1932 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _410_
timestamp 1683767628
transform 1 0 4048 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _411_
timestamp 1683767628
transform 1 0 11684 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _412_
timestamp 1683767628
transform 1 0 5612 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _413_
timestamp 1683767628
transform 1 0 2484 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _414_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1748 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 14168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__CLK
timestamp 1683767628
transform 1 0 13708 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__CLK
timestamp 1683767628
transform 1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__CLK
timestamp 1683767628
transform 1 0 13524 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__CLK
timestamp 1683767628
transform 1 0 8372 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__CLK
timestamp 1683767628
transform 1 0 10672 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__CLK
timestamp 1683767628
transform 1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__CLK
timestamp 1683767628
transform 1 0 12144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__CLK
timestamp 1683767628
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__CLK
timestamp 1683767628
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__CLK
timestamp 1683767628
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__CLK
timestamp 1683767628
transform 1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__CLK
timestamp 1683767628
transform 1 0 11408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__CLK
timestamp 1683767628
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__CLK
timestamp 1683767628
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__CLK
timestamp 1683767628
transform 1 0 13524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__CLK
timestamp 1683767628
transform 1 0 11224 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__CLK
timestamp 1683767628
transform 1 0 13524 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__CLK
timestamp 1683767628
transform 1 0 13800 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__CLK
timestamp 1683767628
transform 1 0 3772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__CLK
timestamp 1683767628
transform 1 0 5980 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__CLK
timestamp 1683767628
transform 1 0 11776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__CLK
timestamp 1683767628
transform 1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__CLK
timestamp 1683767628
transform 1 0 4876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1683767628
transform 1 0 2208 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  fanout1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout2
timestamp 1683767628
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout3
timestamp 1683767628
transform 1 0 10672 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout4
timestamp 1683767628
transform 1 0 14168 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout5
timestamp 1683767628
transform 1 0 11592 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout7
timestamp 1683767628
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout8
timestamp 1683767628
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout9
timestamp 1683767628
transform 1 0 13248 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 16928 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1683767628
transform 1 0 11868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout12
timestamp 1683767628
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1683767628
transform 1 0 12512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp 1683767628
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1683767628
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1683767628
transform 1 0 12144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout17
timestamp 1683767628
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout18
timestamp 1683767628
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout19
timestamp 1683767628
transform 1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1683767628
transform 1 0 4784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1683767628
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1683767628
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout23
timestamp 1683767628
transform 1 0 1840 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 1683767628
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout25
timestamp 1683767628
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1683767628
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1683767628
transform 1 0 11960 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1683767628
transform 1 0 14996 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1683767628
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout30
timestamp 1683767628
transform 1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2116 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2392 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_31
timestamp 1683767628
transform 1 0 3956 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_37
timestamp 1683767628
transform 1 0 4508 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5704 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57
timestamp 1683767628
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_78
timestamp 1683767628
transform 1 0 8280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1683767628
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85
timestamp 1683767628
transform 1 0 8924 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_95
timestamp 1683767628
transform 1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_103
timestamp 1683767628
transform 1 0 10580 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_106
timestamp 1683767628
transform 1 0 10856 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1683767628
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1683767628
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_120 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12144 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_132
timestamp 1683767628
transform 1 0 13248 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_137
timestamp 1683767628
transform 1 0 13708 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1683767628
transform 1 0 14076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_162
timestamp 1683767628
transform 1 0 16008 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1683767628
transform 1 0 16652 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_181 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 17756 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_189
timestamp 1683767628
transform 1 0 18492 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_3
timestamp 1683767628
transform 1 0 1380 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_29
timestamp 1683767628
transform 1 0 3772 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_52
timestamp 1683767628
transform 1 0 5888 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1683767628
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1683767628
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_62
timestamp 1683767628
transform 1 0 6808 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_68
timestamp 1683767628
transform 1 0 7360 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_76
timestamp 1683767628
transform 1 0 8096 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_102
timestamp 1683767628
transform 1 0 10488 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_108
timestamp 1683767628
transform 1 0 11040 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1683767628
transform 1 0 11500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_135
timestamp 1683767628
transform 1 0 13524 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_157
timestamp 1683767628
transform 1 0 15548 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 1683767628
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1683767628
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 1683767628
transform 1 0 17756 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 1683767628
transform 1 0 18492 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 1683767628
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_12
timestamp 1683767628
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_19
timestamp 1683767628
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1683767628
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1683767628
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_33
timestamp 1683767628
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 1683767628
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_52
timestamp 1683767628
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_56
timestamp 1683767628
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_60
timestamp 1683767628
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_66
timestamp 1683767628
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_72
timestamp 1683767628
transform 1 0 7728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_77
timestamp 1683767628
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1683767628
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1683767628
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_90
timestamp 1683767628
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_94
timestamp 1683767628
transform 1 0 9752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_115
timestamp 1683767628
transform 1 0 11684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_120
timestamp 1683767628
transform 1 0 12144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_128
timestamp 1683767628
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_132
timestamp 1683767628
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_136
timestamp 1683767628
transform 1 0 13616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1683767628
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1683767628
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_145
timestamp 1683767628
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_152
timestamp 1683767628
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_163
timestamp 1683767628
transform 1 0 16100 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_175
timestamp 1683767628
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_187
timestamp 1683767628
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_3
timestamp 1683767628
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_9
timestamp 1683767628
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_17
timestamp 1683767628
transform 1 0 2668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_29
timestamp 1683767628
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_36
timestamp 1683767628
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1683767628
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_57
timestamp 1683767628
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_65
timestamp 1683767628
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_72
timestamp 1683767628
transform 1 0 7728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_77
timestamp 1683767628
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_85
timestamp 1683767628
transform 1 0 8924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_96
timestamp 1683767628
transform 1 0 9936 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1683767628
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1683767628
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_135
timestamp 1683767628
transform 1 0 13524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_138
timestamp 1683767628
transform 1 0 13800 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_159
timestamp 1683767628
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_163
timestamp 1683767628
transform 1 0 16100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1683767628
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_169
timestamp 1683767628
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_177
timestamp 1683767628
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_183
timestamp 1683767628
transform 1 0 17940 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_189
timestamp 1683767628
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 1683767628
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_9
timestamp 1683767628
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 1683767628
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1683767628
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1683767628
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 1683767628
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_45
timestamp 1683767628
transform 1 0 5244 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_54
timestamp 1683767628
transform 1 0 6072 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_67
timestamp 1683767628
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1683767628
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1683767628
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1683767628
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_96
timestamp 1683767628
transform 1 0 9936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_119
timestamp 1683767628
transform 1 0 12052 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_122
timestamp 1683767628
transform 1 0 12328 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_133
timestamp 1683767628
transform 1 0 13340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1683767628
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1683767628
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_162
timestamp 1683767628
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_174
timestamp 1683767628
transform 1 0 17112 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_185
timestamp 1683767628
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_189
timestamp 1683767628
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_3
timestamp 1683767628
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_12
timestamp 1683767628
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_35
timestamp 1683767628
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_40
timestamp 1683767628
transform 1 0 4784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_43
timestamp 1683767628
transform 1 0 5060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1683767628
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1683767628
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1683767628
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_62
timestamp 1683767628
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_89
timestamp 1683767628
transform 1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_96
timestamp 1683767628
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_102
timestamp 1683767628
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_107
timestamp 1683767628
transform 1 0 10948 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1683767628
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_113
timestamp 1683767628
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_119
timestamp 1683767628
transform 1 0 12052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_131
timestamp 1683767628
transform 1 0 13156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_137
timestamp 1683767628
transform 1 0 13708 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_158
timestamp 1683767628
transform 1 0 15640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_162
timestamp 1683767628
transform 1 0 16008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 1683767628
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 1683767628
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_179
timestamp 1683767628
transform 1 0 17572 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_187
timestamp 1683767628
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 1683767628
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_11
timestamp 1683767628
transform 1 0 2116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_17
timestamp 1683767628
transform 1 0 2668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1683767628
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_29
timestamp 1683767628
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_33
timestamp 1683767628
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_38
timestamp 1683767628
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_44
timestamp 1683767628
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_48
timestamp 1683767628
transform 1 0 5520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_69
timestamp 1683767628
transform 1 0 7452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_72
timestamp 1683767628
transform 1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1683767628
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1683767628
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1683767628
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_106
timestamp 1683767628
transform 1 0 10856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_109
timestamp 1683767628
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_114
timestamp 1683767628
transform 1 0 11592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_118
timestamp 1683767628
transform 1 0 11960 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_124
timestamp 1683767628
transform 1 0 12512 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_129
timestamp 1683767628
transform 1 0 12972 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_137
timestamp 1683767628
transform 1 0 13708 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1683767628
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_162
timestamp 1683767628
transform 1 0 16008 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_174
timestamp 1683767628
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_186
timestamp 1683767628
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1683767628
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_8
timestamp 1683767628
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_15
timestamp 1683767628
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_21
timestamp 1683767628
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_25
timestamp 1683767628
transform 1 0 3404 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_33
timestamp 1683767628
transform 1 0 4140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_37
timestamp 1683767628
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_43
timestamp 1683767628
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_48
timestamp 1683767628
transform 1 0 5520 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1683767628
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1683767628
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_67
timestamp 1683767628
transform 1 0 7268 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_73
timestamp 1683767628
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_77
timestamp 1683767628
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_82
timestamp 1683767628
transform 1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_87
timestamp 1683767628
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1683767628
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1683767628
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_134
timestamp 1683767628
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_157
timestamp 1683767628
transform 1 0 15548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_161
timestamp 1683767628
transform 1 0 15916 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1683767628
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 1683767628
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_173
timestamp 1683767628
transform 1 0 17020 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_178
timestamp 1683767628
transform 1 0 17480 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1683767628
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_7
timestamp 1683767628
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_11
timestamp 1683767628
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_22
timestamp 1683767628
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1683767628
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_36
timestamp 1683767628
transform 1 0 4416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_45
timestamp 1683767628
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_52
timestamp 1683767628
transform 1 0 5888 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_60
timestamp 1683767628
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1683767628
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_87
timestamp 1683767628
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_92
timestamp 1683767628
transform 1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_97
timestamp 1683767628
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_103
timestamp 1683767628
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_119
timestamp 1683767628
transform 1 0 12052 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_123
timestamp 1683767628
transform 1 0 12420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_129
timestamp 1683767628
transform 1 0 12972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_134
timestamp 1683767628
transform 1 0 13432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1683767628
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 1683767628
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_163
timestamp 1683767628
transform 1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_177
timestamp 1683767628
transform 1 0 17388 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_186
timestamp 1683767628
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_3
timestamp 1683767628
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_7
timestamp 1683767628
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_17
timestamp 1683767628
transform 1 0 2668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_28
timestamp 1683767628
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_38
timestamp 1683767628
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_45
timestamp 1683767628
transform 1 0 5244 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_51
timestamp 1683767628
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1683767628
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1683767628
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_64
timestamp 1683767628
transform 1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_77
timestamp 1683767628
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_81
timestamp 1683767628
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_88
timestamp 1683767628
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_97
timestamp 1683767628
transform 1 0 10028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_104
timestamp 1683767628
transform 1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 1683767628
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1683767628
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_118
timestamp 1683767628
transform 1 0 11960 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_131
timestamp 1683767628
transform 1 0 13156 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_137
timestamp 1683767628
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_140
timestamp 1683767628
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_150
timestamp 1683767628
transform 1 0 14904 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_158
timestamp 1683767628
transform 1 0 15640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1683767628
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp 1683767628
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_175
timestamp 1683767628
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_181
timestamp 1683767628
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 1683767628
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 1683767628
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_11
timestamp 1683767628
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_20
timestamp 1683767628
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1683767628
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_38
timestamp 1683767628
transform 1 0 4600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_50
timestamp 1683767628
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_54
timestamp 1683767628
transform 1 0 6072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_62
timestamp 1683767628
transform 1 0 6808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_77
timestamp 1683767628
transform 1 0 8188 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1683767628
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_85
timestamp 1683767628
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_97
timestamp 1683767628
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_109
timestamp 1683767628
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_118
timestamp 1683767628
transform 1 0 11960 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_130
timestamp 1683767628
transform 1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_136
timestamp 1683767628
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1683767628
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_151
timestamp 1683767628
transform 1 0 14996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_156
timestamp 1683767628
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_170
timestamp 1683767628
transform 1 0 16744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_182
timestamp 1683767628
transform 1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 1683767628
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 1683767628
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_9
timestamp 1683767628
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_19
timestamp 1683767628
transform 1 0 2852 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_26
timestamp 1683767628
transform 1 0 3496 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_38
timestamp 1683767628
transform 1 0 4600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_47
timestamp 1683767628
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 1683767628
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp 1683767628
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_65
timestamp 1683767628
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_76
timestamp 1683767628
transform 1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_86
timestamp 1683767628
transform 1 0 9016 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1683767628
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1683767628
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1683767628
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_122
timestamp 1683767628
transform 1 0 12328 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_128
timestamp 1683767628
transform 1 0 12880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_134
timestamp 1683767628
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_144
timestamp 1683767628
transform 1 0 14352 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_155
timestamp 1683767628
transform 1 0 15364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_164
timestamp 1683767628
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1683767628
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_173
timestamp 1683767628
transform 1 0 17020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_186
timestamp 1683767628
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1683767628
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_9
timestamp 1683767628
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_17
timestamp 1683767628
transform 1 0 2668 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1683767628
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1683767628
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1683767628
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1683767628
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_58
timestamp 1683767628
transform 1 0 6440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_65
timestamp 1683767628
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_72
timestamp 1683767628
transform 1 0 7728 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1683767628
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1683767628
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1683767628
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_104
timestamp 1683767628
transform 1 0 10672 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_113
timestamp 1683767628
transform 1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_122
timestamp 1683767628
transform 1 0 12328 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1683767628
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1683767628
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_149
timestamp 1683767628
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_155
timestamp 1683767628
transform 1 0 15364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_168
timestamp 1683767628
transform 1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_182
timestamp 1683767628
transform 1 0 17848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_187
timestamp 1683767628
transform 1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1683767628
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_9
timestamp 1683767628
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_17
timestamp 1683767628
transform 1 0 2668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_25
timestamp 1683767628
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_34
timestamp 1683767628
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_46
timestamp 1683767628
transform 1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1683767628
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1683767628
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_61
timestamp 1683767628
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_68
timestamp 1683767628
transform 1 0 7360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_75
timestamp 1683767628
transform 1 0 8004 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_81
timestamp 1683767628
transform 1 0 8556 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_85
timestamp 1683767628
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_89
timestamp 1683767628
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_98
timestamp 1683767628
transform 1 0 10120 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 1683767628
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1683767628
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_117
timestamp 1683767628
transform 1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1683767628
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_125
timestamp 1683767628
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_130
timestamp 1683767628
transform 1 0 13064 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_140
timestamp 1683767628
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_145
timestamp 1683767628
transform 1 0 14444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_150
timestamp 1683767628
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_161
timestamp 1683767628
transform 1 0 15916 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1683767628
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 1683767628
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_173
timestamp 1683767628
transform 1 0 17020 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_181
timestamp 1683767628
transform 1 0 17756 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_186
timestamp 1683767628
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1683767628
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_11
timestamp 1683767628
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_16
timestamp 1683767628
transform 1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_20
timestamp 1683767628
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1683767628
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 1683767628
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_37
timestamp 1683767628
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_44
timestamp 1683767628
transform 1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_50
timestamp 1683767628
transform 1 0 5704 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_60
timestamp 1683767628
transform 1 0 6624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_70
timestamp 1683767628
transform 1 0 7544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_76
timestamp 1683767628
transform 1 0 8096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1683767628
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1683767628
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_89
timestamp 1683767628
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_96
timestamp 1683767628
transform 1 0 9936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_101
timestamp 1683767628
transform 1 0 10396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_108
timestamp 1683767628
transform 1 0 11040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_113
timestamp 1683767628
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_121
timestamp 1683767628
transform 1 0 12236 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_126
timestamp 1683767628
transform 1 0 12696 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_131
timestamp 1683767628
transform 1 0 13156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_136
timestamp 1683767628
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1683767628
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_148
timestamp 1683767628
transform 1 0 14720 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_157
timestamp 1683767628
transform 1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_165
timestamp 1683767628
transform 1 0 16284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_172
timestamp 1683767628
transform 1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_181
timestamp 1683767628
transform 1 0 17756 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_186
timestamp 1683767628
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1683767628
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_7
timestamp 1683767628
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_18
timestamp 1683767628
transform 1 0 2760 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_29
timestamp 1683767628
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_41
timestamp 1683767628
transform 1 0 4876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_47
timestamp 1683767628
transform 1 0 5428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1683767628
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_57
timestamp 1683767628
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_70
timestamp 1683767628
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_76
timestamp 1683767628
transform 1 0 8096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_91
timestamp 1683767628
transform 1 0 9476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_98
timestamp 1683767628
transform 1 0 10120 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1683767628
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_113
timestamp 1683767628
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_121
timestamp 1683767628
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_130
timestamp 1683767628
transform 1 0 13064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_139
timestamp 1683767628
transform 1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_151
timestamp 1683767628
transform 1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_157
timestamp 1683767628
transform 1 0 15548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1683767628
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1683767628
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_178
timestamp 1683767628
transform 1 0 17480 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 1683767628
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_11
timestamp 1683767628
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_16
timestamp 1683767628
transform 1 0 2576 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_29
timestamp 1683767628
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_39
timestamp 1683767628
transform 1 0 4692 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_46
timestamp 1683767628
transform 1 0 5336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_53
timestamp 1683767628
transform 1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_61
timestamp 1683767628
transform 1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_75
timestamp 1683767628
transform 1 0 8004 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1683767628
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1683767628
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_93
timestamp 1683767628
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_97
timestamp 1683767628
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_101
timestamp 1683767628
transform 1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_106
timestamp 1683767628
transform 1 0 10856 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_115
timestamp 1683767628
transform 1 0 11684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_122
timestamp 1683767628
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_128
timestamp 1683767628
transform 1 0 12880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1683767628
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1683767628
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_146
timestamp 1683767628
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_150
timestamp 1683767628
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_155
timestamp 1683767628
transform 1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_161
timestamp 1683767628
transform 1 0 15916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_169
timestamp 1683767628
transform 1 0 16652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_175
timestamp 1683767628
transform 1 0 17204 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_187
timestamp 1683767628
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1683767628
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_11
timestamp 1683767628
transform 1 0 2116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_15
timestamp 1683767628
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_24
timestamp 1683767628
transform 1 0 3312 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_43
timestamp 1683767628
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_48
timestamp 1683767628
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1683767628
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_66
timestamp 1683767628
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_74
timestamp 1683767628
transform 1 0 7912 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_90
timestamp 1683767628
transform 1 0 9384 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_99
timestamp 1683767628
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 1683767628
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1683767628
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_123
timestamp 1683767628
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_129
timestamp 1683767628
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_140
timestamp 1683767628
transform 1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_145
timestamp 1683767628
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_157
timestamp 1683767628
transform 1 0 15548 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1683767628
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1683767628
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_176
timestamp 1683767628
transform 1 0 17296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_187
timestamp 1683767628
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1683767628
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_14
timestamp 1683767628
transform 1 0 2392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1683767628
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_29
timestamp 1683767628
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_39
timestamp 1683767628
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_51
timestamp 1683767628
transform 1 0 5796 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_55
timestamp 1683767628
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_59
timestamp 1683767628
transform 1 0 6532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_66
timestamp 1683767628
transform 1 0 7176 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1683767628
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1683767628
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_89
timestamp 1683767628
transform 1 0 9292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_100
timestamp 1683767628
transform 1 0 10304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_111
timestamp 1683767628
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_119
timestamp 1683767628
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_126
timestamp 1683767628
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 1683767628
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1683767628
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_141
timestamp 1683767628
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_145
timestamp 1683767628
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_154
timestamp 1683767628
transform 1 0 15272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_163
timestamp 1683767628
transform 1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_173
timestamp 1683767628
transform 1 0 17020 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_186
timestamp 1683767628
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_3
timestamp 1683767628
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_11
timestamp 1683767628
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_23
timestamp 1683767628
transform 1 0 3220 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_27
timestamp 1683767628
transform 1 0 3588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_33
timestamp 1683767628
transform 1 0 4140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_40
timestamp 1683767628
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_46
timestamp 1683767628
transform 1 0 5336 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1683767628
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1683767628
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_63
timestamp 1683767628
transform 1 0 6900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_69
timestamp 1683767628
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_77
timestamp 1683767628
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_86
timestamp 1683767628
transform 1 0 9016 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_100
timestamp 1683767628
transform 1 0 10304 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1683767628
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1683767628
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_118
timestamp 1683767628
transform 1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_128
timestamp 1683767628
transform 1 0 12880 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_133
timestamp 1683767628
transform 1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_141
timestamp 1683767628
transform 1 0 14076 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_152
timestamp 1683767628
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1683767628
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1683767628
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_178
timestamp 1683767628
transform 1 0 17480 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_3
timestamp 1683767628
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_12
timestamp 1683767628
transform 1 0 2208 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_18
timestamp 1683767628
transform 1 0 2760 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1683767628
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1683767628
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_40
timestamp 1683767628
transform 1 0 4784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_45
timestamp 1683767628
transform 1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_53
timestamp 1683767628
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_61
timestamp 1683767628
transform 1 0 6716 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_74
timestamp 1683767628
transform 1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1683767628
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_85
timestamp 1683767628
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_91
timestamp 1683767628
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_95
timestamp 1683767628
transform 1 0 9844 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_100
timestamp 1683767628
transform 1 0 10304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_111
timestamp 1683767628
transform 1 0 11316 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_119
timestamp 1683767628
transform 1 0 12052 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_123
timestamp 1683767628
transform 1 0 12420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_132
timestamp 1683767628
transform 1 0 13248 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1683767628
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1683767628
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_147
timestamp 1683767628
transform 1 0 14628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_154
timestamp 1683767628
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_163
timestamp 1683767628
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_175
timestamp 1683767628
transform 1 0 17204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_181
timestamp 1683767628
transform 1 0 17756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_189
timestamp 1683767628
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1683767628
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_15
timestamp 1683767628
transform 1 0 2484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_28
timestamp 1683767628
transform 1 0 3680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_37
timestamp 1683767628
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_49
timestamp 1683767628
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1683767628
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 1683767628
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_65
timestamp 1683767628
transform 1 0 7084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_77
timestamp 1683767628
transform 1 0 8188 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_83
timestamp 1683767628
transform 1 0 8740 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_99
timestamp 1683767628
transform 1 0 10212 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 1683767628
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 1683767628
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_121
timestamp 1683767628
transform 1 0 12236 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_134
timestamp 1683767628
transform 1 0 13432 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_146
timestamp 1683767628
transform 1 0 14536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_154
timestamp 1683767628
transform 1 0 15272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_163
timestamp 1683767628
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1683767628
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 1683767628
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_177
timestamp 1683767628
transform 1 0 17388 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_186
timestamp 1683767628
transform 1 0 18216 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1683767628
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1683767628
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1683767628
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 1683767628
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_35
timestamp 1683767628
transform 1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_42
timestamp 1683767628
transform 1 0 4968 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_53
timestamp 1683767628
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_57
timestamp 1683767628
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_65
timestamp 1683767628
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_71
timestamp 1683767628
transform 1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_75
timestamp 1683767628
transform 1 0 8004 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1683767628
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1683767628
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_89
timestamp 1683767628
transform 1 0 9292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_94
timestamp 1683767628
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_103
timestamp 1683767628
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_111
timestamp 1683767628
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_113
timestamp 1683767628
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_117
timestamp 1683767628
transform 1 0 11868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_121
timestamp 1683767628
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_125
timestamp 1683767628
transform 1 0 12604 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_131
timestamp 1683767628
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1683767628
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1683767628
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_149
timestamp 1683767628
transform 1 0 14812 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_155
timestamp 1683767628
transform 1 0 15364 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_160
timestamp 1683767628
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_167
timestamp 1683767628
transform 1 0 16468 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_169
timestamp 1683767628
transform 1 0 16652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_177
timestamp 1683767628
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_182
timestamp 1683767628
transform 1 0 17848 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1683767628
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1683767628
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1683767628
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1683767628
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1683767628
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1683767628
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1683767628
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1683767628
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1683767628
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1683767628
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1683767628
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1683767628
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1683767628
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1683767628
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1683767628
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1683767628
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1683767628
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1683767628
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1683767628
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1683767628
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1683767628
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1683767628
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1683767628
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1683767628
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1683767628
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1683767628
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1683767628
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1683767628
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1683767628
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1683767628
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1683767628
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1683767628
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1683767628
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1683767628
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1683767628
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1683767628
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1683767628
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1683767628
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1683767628
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1683767628
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1683767628
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1683767628
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1683767628
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1683767628
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1683767628
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1683767628
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1683767628
transform 1 0 6256 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 6440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5704 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3588 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[0\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5980 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[0\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1683767628
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1683767628
transform 1 0 5704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1683767628
transform 1 0 3864 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1683767628
transform 1 0 4876 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1683767628
transform 1 0 3128 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[1\].id.delayenb1
timestamp 1683767628
transform 1 0 5520 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1683767628
transform 1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1683767628
transform 1 0 4324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1683767628
transform 1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1683767628
transform 1 0 14168 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1683767628
transform 1 0 14168 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1683767628
transform 1 0 14628 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[2\].id.delayenb1
timestamp 1683767628
transform 1 0 13616 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1683767628
transform 1 0 14996 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1683767628
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1683767628
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1683767628
transform 1 0 11592 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1683767628
transform 1 0 12696 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1683767628
transform 1 0 10672 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[3\].id.delayenb1
timestamp 1683767628
transform 1 0 12972 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1683767628
transform 1 0 11960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1683767628
transform 1 0 7268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1683767628
transform 1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1683767628
transform 1 0 4416 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1683767628
transform 1 0 6256 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp 1683767628
transform 1 0 4048 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[4\].id.delayenb1
timestamp 1683767628
transform 1 0 6992 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1683767628
transform 1 0 5888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1683767628
transform 1 0 4968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1683767628
transform 1 0 3312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1683767628
transform 1 0 1748 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1683767628
transform 1 0 2852 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb0
timestamp 1683767628
transform 1 0 1472 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1683767628
transform 1 0 2944 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1683767628
transform 1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1683767628
transform 1 0 2392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1683767628
transform 1 0 4692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1683767628
transform 1 0 4140 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1683767628
transform 1 0 3864 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1683767628
transform 1 0 3864 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1683767628
transform 1 0 3036 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1683767628
transform 1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1683767628
transform 1 0 5704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1683767628
transform 1 0 9016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1683767628
transform 1 0 7268 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1683767628
transform 1 0 8096 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1683767628
transform 1 0 6440 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[7\].id.delayenb1
timestamp 1683767628
transform 1 0 8280 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1683767628
transform 1 0 9476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1683767628
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1683767628
transform 1 0 17572 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1683767628
transform 1 0 16744 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1683767628
transform 1 0 17296 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1683767628
transform 1 0 15456 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1683767628
transform 1 0 16744 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1683767628
transform 1 0 16192 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1683767628
transform 1 0 18124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1683767628
transform 1 0 16192 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1683767628
transform 1 0 17664 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1683767628
transform 1 0 17756 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp 1683767628
transform 1 0 16836 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1683767628
transform 1 0 16376 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1683767628
transform 1 0 17940 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1683767628
transform 1 0 17940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1683767628
transform 1 0 16652 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1683767628
transform 1 0 17112 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1683767628
transform 1 0 16836 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1683767628
transform 1 0 16836 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[10\].id.delayenb1
timestamp 1683767628
transform 1 0 16744 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1683767628
transform 1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1683767628
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1683767628
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 17204 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1
timestamp 1683767628
transform 1 0 18032 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 16836 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[11\].id.delayenb1
timestamp 1683767628
transform 1 0 17296 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1683767628
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 11592 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10856 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10
timestamp 1683767628
transform 1 0 2300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  ringosc.ibufp11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2024 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 17204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 15732 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1683767628
transform 1 0 16744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1683767628
transform 1 0 15548 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1683767628
transform 1 0 15824 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1683767628
transform 1 0 15732 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_1  ringosc.iss.delayenb1
timestamp 1683767628
transform 1 0 15456 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.iss.delayint0
timestamp 1683767628
transform 1 0 16744 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1683767628
transform 1 0 16376 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1683767628
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1683767628
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1683767628
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1683767628
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1683767628
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1683767628
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1683767628
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1683767628
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1683767628
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1683767628
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1683767628
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1683767628
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1683767628
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1683767628
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1683767628
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1683767628
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1683767628
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1683767628
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1683767628
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1683767628
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1683767628
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1683767628
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1683767628
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1683767628
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1683767628
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1683767628
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1683767628
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1683767628
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1683767628
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1683767628
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1683767628
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1683767628
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1683767628
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1683767628
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1683767628
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1683767628
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1683767628
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1683767628
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1683767628
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1683767628
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1683767628
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1683767628
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1683767628
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1683767628
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1683767628
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1683767628
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1683767628
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1683767628
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1683767628
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1683767628
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1683767628
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1683767628
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1683767628
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1683767628
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1683767628
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1683767628
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1683767628
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1683767628
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1683767628
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1683767628
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1683767628
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1683767628
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1683767628
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1683767628
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1683767628
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1683767628
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1683767628
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1683767628
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1683767628
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1683767628
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1683767628
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1683767628
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1683767628
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1683767628
transform 1 0 16560 0 1 13056
box -38 -48 130 592
<< labels >>
flabel metal4 s 8208 1040 8528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16208 1040 16528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 1040 4528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12208 1040 12528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 5538 14200 5594 15000 0 FreeSans 224 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 7010 14200 7066 15000 0 FreeSans 224 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 8482 14200 8538 15000 0 FreeSans 224 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 9954 14200 10010 15000 0 FreeSans 224 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 11426 14200 11482 15000 0 FreeSans 224 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 12898 14200 12954 15000 0 FreeSans 224 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 14370 14200 14426 15000 0 FreeSans 224 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 15842 14200 15898 15000 0 FreeSans 224 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 17314 14200 17370 15000 0 FreeSans 224 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 18786 14200 18842 15000 0 FreeSans 224 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 19200 13336 20000 13456 0 FreeSans 480 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 19200 10888 20000 11008 0 FreeSans 480 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 19200 8440 20000 8560 0 FreeSans 480 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 19200 5992 20000 6112 0 FreeSans 480 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 19200 3544 20000 3664 0 FreeSans 480 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 19200 1096 20000 1216 0 FreeSans 480 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 1122 14200 1178 15000 0 FreeSans 224 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 2594 14200 2650 15000 0 FreeSans 224 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 4066 14200 4122 15000 0 FreeSans 224 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 resetb
port 38 nsew signal input
rlabel metal1 9982 13056 9982 13056 0 VGND
rlabel metal1 9982 13600 9982 13600 0 VPWR
rlabel metal1 15877 3094 15877 3094 0 _000_
rlabel metal1 13386 3434 13386 3434 0 _001_
rlabel metal1 16238 4148 16238 4148 0 _002_
rlabel metal2 7038 1768 7038 1768 0 _003_
rlabel metal1 10810 1462 10810 1462 0 _004_
rlabel metal2 10902 2210 10902 2210 0 _005_
rlabel metal1 11737 3434 11737 3434 0 _006_
rlabel metal1 7176 4250 7176 4250 0 _007_
rlabel metal1 9108 4998 9108 4998 0 _008_
rlabel metal1 8096 5338 8096 5338 0 _009_
rlabel metal1 9883 5270 9883 5270 0 _010_
rlabel metal2 12650 5032 12650 5032 0 _011_
rlabel metal1 15877 4522 15877 4522 0 _012_
rlabel metal2 16882 5474 16882 5474 0 _013_
rlabel metal1 14299 5270 14299 5270 0 _014_
rlabel metal2 11914 1734 11914 1734 0 _015_
rlabel metal1 14391 2006 14391 2006 0 _016_
rlabel metal2 14950 1768 14950 1768 0 _017_
rlabel metal1 3733 2006 3733 2006 0 _018_
rlabel metal1 4554 1530 4554 1530 0 _019_
rlabel metal2 13018 2856 13018 2856 0 _020_
rlabel metal1 7038 4631 7038 4631 0 _021_
rlabel metal1 4646 4148 4646 4148 0 _022_
rlabel metal1 15778 2958 15778 2958 0 _023_
rlabel metal1 17342 3604 17342 3604 0 _024_
rlabel metal1 15456 4046 15456 4046 0 _025_
rlabel metal1 6660 1530 6660 1530 0 _026_
rlabel metal1 9108 1530 9108 1530 0 _027_
rlabel metal1 10350 1462 10350 1462 0 _028_
rlabel metal1 9844 3434 9844 3434 0 _029_
rlabel metal1 7590 3706 7590 3706 0 _030_
rlabel metal1 9016 4658 9016 4658 0 _031_
rlabel metal2 7130 5916 7130 5916 0 _032_
rlabel metal1 9476 5270 9476 5270 0 _033_
rlabel metal2 11914 6256 11914 6256 0 _034_
rlabel metal1 14444 4522 14444 4522 0 _035_
rlabel metal2 14490 6188 14490 6188 0 _036_
rlabel metal2 14030 5712 14030 5712 0 _037_
rlabel metal2 2622 1666 2622 1666 0 _038_
rlabel metal2 4922 1700 4922 1700 0 _039_
rlabel metal1 11592 2958 11592 2958 0 _040_
rlabel metal1 6210 4658 6210 4658 0 _041_
rlabel metal2 2806 4318 2806 4318 0 _042_
rlabel metal1 7912 3162 7912 3162 0 _043_
rlabel metal2 10718 9282 10718 9282 0 _044_
rlabel metal1 8234 7242 8234 7242 0 _045_
rlabel metal1 13846 10642 13846 10642 0 _046_
rlabel metal1 9200 8262 9200 8262 0 _047_
rlabel metal1 2300 5678 2300 5678 0 _048_
rlabel metal1 2070 5270 2070 5270 0 _049_
rlabel via1 1886 2414 1886 2414 0 _050_
rlabel metal1 15134 2550 15134 2550 0 _051_
rlabel metal1 2806 7344 2806 7344 0 _052_
rlabel metal2 5014 7174 5014 7174 0 _053_
rlabel metal2 5474 5882 5474 5882 0 _054_
rlabel metal1 5198 5338 5198 5338 0 _055_
rlabel metal1 5612 5746 5612 5746 0 _056_
rlabel metal2 6026 5508 6026 5508 0 _057_
rlabel metal1 6578 2448 6578 2448 0 _058_
rlabel metal1 4922 5168 4922 5168 0 _059_
rlabel metal1 6164 2414 6164 2414 0 _060_
rlabel metal1 5934 2618 5934 2618 0 _061_
rlabel metal1 4945 3502 4945 3502 0 _062_
rlabel metal1 3404 2618 3404 2618 0 _063_
rlabel metal1 4784 2414 4784 2414 0 _064_
rlabel metal1 4876 2618 4876 2618 0 _065_
rlabel metal1 5060 5202 5060 5202 0 _066_
rlabel metal1 4876 7310 4876 7310 0 _067_
rlabel metal1 2668 7378 2668 7378 0 _068_
rlabel metal1 3266 7310 3266 7310 0 _069_
rlabel metal1 2392 7174 2392 7174 0 _070_
rlabel metal1 5934 4046 5934 4046 0 _071_
rlabel metal1 2254 5168 2254 5168 0 _072_
rlabel metal2 4738 5406 4738 5406 0 _073_
rlabel metal1 2714 5644 2714 5644 0 _074_
rlabel metal1 3174 5168 3174 5168 0 _075_
rlabel metal2 3358 6188 3358 6188 0 _076_
rlabel metal2 2438 6120 2438 6120 0 _077_
rlabel metal2 2254 6222 2254 6222 0 _078_
rlabel metal2 2530 6596 2530 6596 0 _079_
rlabel metal1 1932 4590 1932 4590 0 _080_
rlabel metal2 1886 4284 1886 4284 0 _081_
rlabel metal1 2254 3502 2254 3502 0 _082_
rlabel metal1 2392 2618 2392 2618 0 _083_
rlabel metal1 2346 3060 2346 3060 0 _084_
rlabel metal1 2438 3570 2438 3570 0 _085_
rlabel metal1 1748 4114 1748 4114 0 _086_
rlabel metal1 2070 6426 2070 6426 0 _087_
rlabel metal1 2714 7208 2714 7208 0 _088_
rlabel metal1 2438 7820 2438 7820 0 _089_
rlabel metal1 6762 7820 6762 7820 0 _090_
rlabel metal1 10810 9894 10810 9894 0 _091_
rlabel metal2 13570 9044 13570 9044 0 _092_
rlabel metal2 14214 8772 14214 8772 0 _093_
rlabel metal2 12926 9316 12926 9316 0 _094_
rlabel metal1 12466 8840 12466 8840 0 _095_
rlabel metal1 10350 9078 10350 9078 0 _096_
rlabel metal2 7130 8126 7130 8126 0 _097_
rlabel metal2 8142 7684 8142 7684 0 _098_
rlabel metal1 10902 6426 10902 6426 0 _099_
rlabel metal1 7314 6902 7314 6902 0 _100_
rlabel metal2 17066 5338 17066 5338 0 _101_
rlabel metal2 3726 3298 3726 3298 0 _102_
rlabel metal1 2852 3706 2852 3706 0 _103_
rlabel metal1 7452 6698 7452 6698 0 _104_
rlabel metal2 8142 7140 8142 7140 0 _105_
rlabel metal1 10258 6426 10258 6426 0 _106_
rlabel metal1 7728 9418 7728 9418 0 _107_
rlabel metal1 11638 11730 11638 11730 0 _108_
rlabel metal2 7866 7548 7866 7548 0 _109_
rlabel metal2 8510 6970 8510 6970 0 _110_
rlabel metal1 13478 7888 13478 7888 0 _111_
rlabel metal1 14260 8262 14260 8262 0 _112_
rlabel metal1 13524 8466 13524 8466 0 _113_
rlabel metal1 14536 7854 14536 7854 0 _114_
rlabel metal1 8970 10676 8970 10676 0 _115_
rlabel metal2 10258 7684 10258 7684 0 _116_
rlabel metal1 10396 7922 10396 7922 0 _117_
rlabel metal2 13294 8228 13294 8228 0 _118_
rlabel metal2 12742 7242 12742 7242 0 _119_
rlabel metal1 12880 6766 12880 6766 0 _120_
rlabel metal1 12834 5882 12834 5882 0 _121_
rlabel metal2 12834 6460 12834 6460 0 _122_
rlabel metal2 13846 7820 13846 7820 0 _123_
rlabel metal1 14490 6834 14490 6834 0 _124_
rlabel metal1 14674 6426 14674 6426 0 _125_
rlabel metal1 10350 6664 10350 6664 0 _126_
rlabel metal1 11040 7310 11040 7310 0 _127_
rlabel metal1 9614 6630 9614 6630 0 _128_
rlabel metal1 6486 6800 6486 6800 0 _129_
rlabel metal1 7314 6426 7314 6426 0 _130_
rlabel metal1 8924 5338 8924 5338 0 _131_
rlabel metal2 9614 3808 9614 3808 0 _132_
rlabel metal1 8970 3910 8970 3910 0 _133_
rlabel metal2 9706 3332 9706 3332 0 _134_
rlabel metal2 6578 2142 6578 2142 0 _135_
rlabel metal1 8510 2550 8510 2550 0 _136_
rlabel metal1 10350 1292 10350 1292 0 _137_
rlabel metal2 9798 1530 9798 1530 0 _138_
rlabel metal2 2990 8364 2990 8364 0 _139_
rlabel metal2 7682 8636 7682 8636 0 _140_
rlabel metal2 9246 10761 9246 10761 0 _141_
rlabel metal2 13570 11084 13570 11084 0 _142_
rlabel metal1 14766 9078 14766 9078 0 _143_
rlabel metal2 9982 10166 9982 10166 0 _144_
rlabel metal2 8510 11322 8510 11322 0 _145_
rlabel metal1 9614 11254 9614 11254 0 _146_
rlabel metal1 8694 11798 8694 11798 0 _147_
rlabel metal1 12650 11016 12650 11016 0 _148_
rlabel metal1 14858 9520 14858 9520 0 _149_
rlabel metal2 15134 8398 15134 8398 0 _150_
rlabel metal1 6624 12410 6624 12410 0 _151_
rlabel metal1 7866 11764 7866 11764 0 _152_
rlabel metal2 15502 10982 15502 10982 0 _153_
rlabel metal2 10258 12274 10258 12274 0 _154_
rlabel metal1 10672 11730 10672 11730 0 _155_
rlabel metal1 13156 10234 13156 10234 0 _156_
rlabel metal1 6716 11322 6716 11322 0 _157_
rlabel metal1 10488 10778 10488 10778 0 _158_
rlabel metal1 6624 13226 6624 13226 0 _159_
rlabel metal1 9016 11186 9016 11186 0 _160_
rlabel metal1 6394 10064 6394 10064 0 _161_
rlabel metal1 7682 9350 7682 9350 0 _162_
rlabel metal1 7682 9622 7682 9622 0 _163_
rlabel metal1 13432 9554 13432 9554 0 _164_
rlabel metal1 14950 11152 14950 11152 0 _165_
rlabel metal2 7498 10132 7498 10132 0 _166_
rlabel metal1 12972 11798 12972 11798 0 _167_
rlabel metal2 12650 11696 12650 11696 0 _168_
rlabel metal1 9200 10234 9200 10234 0 _169_
rlabel metal1 9246 10778 9246 10778 0 _170_
rlabel metal1 9568 11186 9568 11186 0 _171_
rlabel metal2 12098 11186 12098 11186 0 _172_
rlabel metal2 13110 10336 13110 10336 0 _173_
rlabel metal1 14490 13158 14490 13158 0 _174_
rlabel metal1 14398 9418 14398 9418 0 _175_
rlabel metal1 14858 11016 14858 11016 0 _176_
rlabel metal2 14766 10948 14766 10948 0 _177_
rlabel metal2 10166 9180 10166 9180 0 _178_
rlabel metal1 9982 9078 9982 9078 0 _179_
rlabel metal1 13754 9350 13754 9350 0 _180_
rlabel metal2 15042 10404 15042 10404 0 _181_
rlabel metal3 866 1156 866 1156 0 clockp[0]
rlabel metal3 2108 1972 2108 1972 0 clockp[1]
rlabel metal2 10166 7072 10166 7072 0 dco
rlabel metal1 2254 2992 2254 2992 0 div[0]
rlabel metal1 1518 3502 1518 3502 0 div[1]
rlabel metal3 820 4420 820 4420 0 div[2]
rlabel metal2 1886 5457 1886 5457 0 div[3]
rlabel metal2 2438 7174 2438 7174 0 div[4]
rlabel metal1 6440 2074 6440 2074 0 dll_control.clock
rlabel metal1 8188 1530 8188 1530 0 dll_control.count0\[0\]
rlabel metal1 5474 2380 5474 2380 0 dll_control.count0\[1\]
rlabel metal1 11454 2618 11454 2618 0 dll_control.count0\[2\]
rlabel metal1 9522 3536 9522 3536 0 dll_control.count0\[3\]
rlabel metal1 2024 7378 2024 7378 0 dll_control.count0\[4\]
rlabel metal1 3266 2448 3266 2448 0 dll_control.count1\[0\]
rlabel metal1 5612 2414 5612 2414 0 dll_control.count1\[1\]
rlabel metal1 10994 3128 10994 3128 0 dll_control.count1\[2\]
rlabel metal1 6808 5134 6808 5134 0 dll_control.count1\[3\]
rlabel metal2 1702 7140 1702 7140 0 dll_control.count1\[4\]
rlabel metal1 14030 2040 14030 2040 0 dll_control.oscbuf\[0\]
rlabel metal2 15502 1564 15502 1564 0 dll_control.oscbuf\[1\]
rlabel metal2 15778 2006 15778 2006 0 dll_control.oscbuf\[2\]
rlabel metal1 16974 3094 16974 3094 0 dll_control.prep\[0\]
rlabel viali 16894 3502 16894 3502 0 dll_control.prep\[1\]
rlabel metal1 17250 3978 17250 3978 0 dll_control.prep\[2\]
rlabel metal1 10902 6630 10902 6630 0 dll_control.tint\[0\]
rlabel metal2 13202 6562 13202 6562 0 dll_control.tint\[1\]
rlabel metal2 15226 7565 15226 7565 0 dll_control.tint\[2\]
rlabel metal2 14582 6188 14582 6188 0 dll_control.tint\[3\]
rlabel metal2 15502 6018 15502 6018 0 dll_control.tint\[4\]
rlabel metal1 9844 5678 9844 5678 0 dll_control.tval\[0\]
rlabel metal2 8602 6086 8602 6086 0 dll_control.tval\[1\]
rlabel metal2 4002 6477 4002 6477 0 enable
rlabel metal3 958 8500 958 8500 0 ext_trim[0]
rlabel metal2 5566 13814 5566 13814 0 ext_trim[10]
rlabel viali 8385 11118 8385 11118 0 ext_trim[11]
rlabel metal2 8563 14348 8563 14348 0 ext_trim[12]
rlabel metal2 10028 11220 10028 11220 0 ext_trim[13]
rlabel metal2 11454 12505 11454 12505 0 ext_trim[14]
rlabel viali 12650 11729 12650 11729 0 ext_trim[15]
rlabel metal1 16054 12852 16054 12852 0 ext_trim[16]
rlabel metal1 15479 11050 15479 11050 0 ext_trim[17]
rlabel metal2 17342 13377 17342 13377 0 ext_trim[18]
rlabel metal1 13294 12206 13294 12206 0 ext_trim[19]
rlabel metal3 1004 9316 1004 9316 0 ext_trim[1]
rlabel metal1 10097 12886 10097 12886 0 ext_trim[20]
rlabel metal1 16192 11118 16192 11118 0 ext_trim[21]
rlabel metal3 17488 8500 17488 8500 0 ext_trim[22]
rlabel metal1 16330 9520 16330 9520 0 ext_trim[23]
rlabel metal1 16146 6256 16146 6256 0 ext_trim[24]
rlabel metal3 17940 1224 17940 1224 0 ext_trim[25]
rlabel metal2 14214 9877 14214 9877 0 ext_trim[2]
rlabel metal3 2499 10948 2499 10948 0 ext_trim[3]
rlabel via2 3726 11781 3726 11781 0 ext_trim[4]
rlabel metal3 1418 12580 1418 12580 0 ext_trim[5]
rlabel metal3 2108 13396 2108 13396 0 ext_trim[6]
rlabel via1 1426 14331 1426 14331 0 ext_trim[7]
rlabel metal2 2622 12505 2622 12505 0 ext_trim[8]
rlabel metal2 4041 14348 4041 14348 0 ext_trim[9]
rlabel metal1 8050 6188 8050 6188 0 net1
rlabel metal2 15778 6460 15778 6460 0 net10
rlabel metal1 7544 9962 7544 9962 0 net11
rlabel metal1 14582 6358 14582 6358 0 net12
rlabel metal2 8878 10642 8878 10642 0 net13
rlabel metal2 4094 2074 4094 2074 0 net14
rlabel metal2 5244 1258 5244 1258 0 net15
rlabel metal2 10810 1632 10810 1632 0 net16
rlabel metal1 14858 2448 14858 2448 0 net17
rlabel metal1 16744 5202 16744 5202 0 net18
rlabel metal1 7958 4522 7958 4522 0 net19
rlabel metal1 12834 8398 12834 8398 0 net2
rlabel metal1 4554 1326 4554 1326 0 net20
rlabel metal1 7084 13158 7084 13158 0 net21
rlabel metal1 2116 12070 2116 12070 0 net22
rlabel metal1 5014 4590 5014 4590 0 net23
rlabel metal1 14996 2414 14996 2414 0 net24
rlabel metal1 16192 5202 16192 5202 0 net25
rlabel metal1 11316 1938 11316 1938 0 net26
rlabel metal1 12282 10608 12282 10608 0 net27
rlabel metal1 14674 9588 14674 9588 0 net28
rlabel metal1 15088 7854 15088 7854 0 net29
rlabel metal2 10718 8398 10718 8398 0 net3
rlabel metal2 13018 6545 13018 6545 0 net30
rlabel metal1 7314 8500 7314 8500 0 net4
rlabel metal1 9752 8942 9752 8942 0 net5
rlabel metal1 13570 10574 13570 10574 0 net6
rlabel metal1 9936 3502 9936 3502 0 net7
rlabel metal1 16238 3502 16238 3502 0 net8
rlabel metal1 10396 8942 10396 8942 0 net9
rlabel metal2 14950 823 14950 823 0 osc
rlabel metal2 4968 4556 4968 4556 0 resetb
rlabel metal2 11822 5882 11822 5882 0 ringosc.c\[0\]
rlabel metal1 2277 9894 2277 9894 0 ringosc.c\[1\]
rlabel metal1 6302 8330 6302 8330 0 ringosc.dstage\[0\].id.d0
rlabel metal2 6118 8772 6118 8772 0 ringosc.dstage\[0\].id.d1
rlabel metal1 5198 7922 5198 7922 0 ringosc.dstage\[0\].id.d2
rlabel metal1 8464 8330 8464 8330 0 ringosc.dstage\[0\].id.in
rlabel metal1 4830 7990 4830 7990 0 ringosc.dstage\[0\].id.out
rlabel metal1 3542 8058 3542 8058 0 ringosc.dstage\[0\].id.trim\[0\]
rlabel metal1 5980 8466 5980 8466 0 ringosc.dstage\[0\].id.trim\[1\]
rlabel metal1 6670 8500 6670 8500 0 ringosc.dstage\[0\].id.ts
rlabel metal1 16974 9146 16974 9146 0 ringosc.dstage\[10\].id.d0
rlabel metal1 17572 10166 17572 10166 0 ringosc.dstage\[10\].id.d1
rlabel metal1 17917 8874 17917 8874 0 ringosc.dstage\[10\].id.d2
rlabel metal2 18170 11118 18170 11118 0 ringosc.dstage\[10\].id.in
rlabel metal2 17618 9214 17618 9214 0 ringosc.dstage\[10\].id.out
rlabel via2 17158 8925 17158 8925 0 ringosc.dstage\[10\].id.trim\[0\]
rlabel metal2 16790 9826 16790 9826 0 ringosc.dstage\[10\].id.trim\[1\]
rlabel metal1 17710 9962 17710 9962 0 ringosc.dstage\[10\].id.ts
rlabel metal1 18216 5882 18216 5882 0 ringosc.dstage\[11\].id.d0
rlabel metal1 18400 6630 18400 6630 0 ringosc.dstage\[11\].id.d1
rlabel metal2 18170 7548 18170 7548 0 ringosc.dstage\[11\].id.d2
rlabel metal2 16974 7990 16974 7990 0 ringosc.dstage\[11\].id.out
rlabel metal1 17066 7310 17066 7310 0 ringosc.dstage\[11\].id.trim\[0\]
rlabel metal2 17342 6528 17342 6528 0 ringosc.dstage\[11\].id.trim\[1\]
rlabel metal2 17802 8092 17802 8092 0 ringosc.dstage\[11\].id.ts
rlabel metal1 5520 10166 5520 10166 0 ringosc.dstage\[1\].id.d0
rlabel metal1 5612 9894 5612 9894 0 ringosc.dstage\[1\].id.d1
rlabel metal1 4600 9010 4600 9010 0 ringosc.dstage\[1\].id.d2
rlabel metal1 4508 9078 4508 9078 0 ringosc.dstage\[1\].id.out
rlabel metal2 3082 9350 3082 9350 0 ringosc.dstage\[1\].id.trim\[0\]
rlabel metal2 5566 9996 5566 9996 0 ringosc.dstage\[1\].id.trim\[1\]
rlabel metal2 5014 9350 5014 9350 0 ringosc.dstage\[1\].id.ts
rlabel metal2 14858 12036 14858 12036 0 ringosc.dstage\[2\].id.d0
rlabel metal2 14582 11968 14582 11968 0 ringosc.dstage\[2\].id.d1
rlabel metal1 14973 12410 14973 12410 0 ringosc.dstage\[2\].id.d2
rlabel via1 14582 12750 14582 12750 0 ringosc.dstage\[2\].id.out
rlabel metal1 14582 12818 14582 12818 0 ringosc.dstage\[2\].id.trim\[0\]
rlabel metal1 13938 11730 13938 11730 0 ringosc.dstage\[2\].id.trim\[1\]
rlabel metal1 8602 10132 8602 10132 0 ringosc.dstage\[2\].id.ts
rlabel metal1 13248 13430 13248 13430 0 ringosc.dstage\[3\].id.d0
rlabel metal1 12880 13158 12880 13158 0 ringosc.dstage\[3\].id.d1
rlabel metal2 12190 13022 12190 13022 0 ringosc.dstage\[3\].id.d2
rlabel metal1 12098 12920 12098 12920 0 ringosc.dstage\[3\].id.out
rlabel metal1 10948 12206 10948 12206 0 ringosc.dstage\[3\].id.trim\[0\]
rlabel metal1 13018 12716 13018 12716 0 ringosc.dstage\[3\].id.trim\[1\]
rlabel metal1 13524 13294 13524 13294 0 ringosc.dstage\[3\].id.ts
rlabel metal1 6302 11866 6302 11866 0 ringosc.dstage\[4\].id.d0
rlabel metal1 6624 12070 6624 12070 0 ringosc.dstage\[4\].id.d1
rlabel metal1 5290 10710 5290 10710 0 ringosc.dstage\[4\].id.d2
rlabel metal1 4876 11322 4876 11322 0 ringosc.dstage\[4\].id.out
rlabel metal2 4094 11322 4094 11322 0 ringosc.dstage\[4\].id.trim\[0\]
rlabel metal1 13846 11186 13846 11186 0 ringosc.dstage\[4\].id.trim\[1\]
rlabel metal1 5980 11730 5980 11730 0 ringosc.dstage\[4\].id.ts
rlabel metal1 3312 10642 3312 10642 0 ringosc.dstage\[5\].id.d0
rlabel metal1 2540 10642 2540 10642 0 ringosc.dstage\[5\].id.d1
rlabel via1 2369 10778 2369 10778 0 ringosc.dstage\[5\].id.d2
rlabel metal2 2254 10540 2254 10540 0 ringosc.dstage\[5\].id.out
rlabel metal2 1518 11900 1518 11900 0 ringosc.dstage\[5\].id.trim\[0\]
rlabel metal2 10626 10336 10626 10336 0 ringosc.dstage\[5\].id.trim\[1\]
rlabel metal1 3588 11730 3588 11730 0 ringosc.dstage\[5\].id.ts
rlabel metal1 4508 13430 4508 13430 0 ringosc.dstage\[6\].id.d0
rlabel metal1 4554 13158 4554 13158 0 ringosc.dstage\[6\].id.d1
rlabel metal1 4945 12138 4945 12138 0 ringosc.dstage\[6\].id.d2
rlabel metal1 5106 12886 5106 12886 0 ringosc.dstage\[6\].id.out
rlabel metal1 3634 12274 3634 12274 0 ringosc.dstage\[6\].id.trim\[0\]
rlabel metal2 13202 12682 13202 12682 0 ringosc.dstage\[6\].id.trim\[1\]
rlabel metal1 4462 12784 4462 12784 0 ringosc.dstage\[6\].id.ts
rlabel metal1 8786 13430 8786 13430 0 ringosc.dstage\[7\].id.d0
rlabel metal1 8924 13158 8924 13158 0 ringosc.dstage\[7\].id.d1
rlabel metal1 8763 13362 8763 13362 0 ringosc.dstage\[7\].id.d2
rlabel metal1 15594 13328 15594 13328 0 ringosc.dstage\[7\].id.out
rlabel metal1 6716 12818 6716 12818 0 ringosc.dstage\[7\].id.trim\[0\]
rlabel metal1 8924 12818 8924 12818 0 ringosc.dstage\[7\].id.trim\[1\]
rlabel metal1 7038 12784 7038 12784 0 ringosc.dstage\[7\].id.ts
rlabel metal1 17664 12274 17664 12274 0 ringosc.dstage\[8\].id.d0
rlabel metal1 16974 12886 16974 12886 0 ringosc.dstage\[8\].id.d1
rlabel metal1 16951 13362 16951 13362 0 ringosc.dstage\[8\].id.d2
rlabel metal1 17342 13226 17342 13226 0 ringosc.dstage\[8\].id.out
rlabel metal2 16790 13124 16790 13124 0 ringosc.dstage\[8\].id.trim\[0\]
rlabel metal2 17342 11764 17342 11764 0 ringosc.dstage\[8\].id.trim\[1\]
rlabel metal1 17342 12784 17342 12784 0 ringosc.dstage\[8\].id.ts
rlabel metal1 17204 11254 17204 11254 0 ringosc.dstage\[9\].id.d0
rlabel via1 18065 12818 18065 12818 0 ringosc.dstage\[9\].id.d1
rlabel metal1 18193 12614 18193 12614 0 ringosc.dstage\[9\].id.d2
rlabel metal1 16882 11764 16882 11764 0 ringosc.dstage\[9\].id.trim\[0\]
rlabel metal1 16422 11084 16422 11084 0 ringosc.dstage\[9\].id.trim\[1\]
rlabel metal2 17434 11900 17434 11900 0 ringosc.dstage\[9\].id.ts
rlabel metal2 15778 6970 15778 6970 0 ringosc.iss.ctrl0
rlabel metal2 16790 8228 16790 8228 0 ringosc.iss.d0
rlabel metal1 16054 8806 16054 8806 0 ringosc.iss.d1
rlabel metal1 16560 7854 16560 7854 0 ringosc.iss.d2
rlabel metal2 17250 5508 17250 5508 0 ringosc.iss.one
rlabel metal1 4462 5202 4462 5202 0 ringosc.iss.reset
rlabel metal1 15824 7922 15824 7922 0 ringosc.iss.trim\[0\]
rlabel metal1 15686 9078 15686 9078 0 ringosc.iss.trim\[1\]
<< properties >>
string FIXED_BBOX 0 0 20000 15000
<< end >>
