VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO picosoc
  CLASS BLOCK ;
  FOREIGN picosoc ;
  ORIGIN 0.000 0.000 ;
  SIZE 2200.000 BY 1500.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.070 10.640 17.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 10.640 57.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.070 10.640 97.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.070 1046.620 97.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.070 10.640 137.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.070 1046.620 137.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.070 10.640 177.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.070 1046.620 177.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.070 10.640 217.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.070 1046.620 217.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.070 10.640 257.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.070 1047.240 257.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.070 10.640 297.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.070 1046.620 297.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.070 10.640 337.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.070 1046.620 337.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.070 10.640 377.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.070 1046.620 377.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.070 10.640 417.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.070 1046.620 417.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.070 10.640 457.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.070 1047.240 457.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 494.070 10.640 497.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 494.070 1046.620 497.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.070 10.640 537.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.070 1046.620 537.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.070 10.640 577.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.070 1046.620 577.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.070 10.640 617.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.070 1047.240 617.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.070 10.640 657.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.070 1046.620 657.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.070 10.640 697.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.070 1046.620 697.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 734.070 10.640 737.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 734.070 1046.620 737.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 774.070 10.640 777.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 774.070 1046.620 777.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.070 10.640 817.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.070 10.640 857.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.070 10.640 897.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 934.070 10.640 937.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.070 10.640 977.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1014.070 10.640 1017.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.070 10.640 1057.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1094.070 10.640 1097.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1134.070 10.640 1137.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1174.070 10.640 1177.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1214.070 10.640 1217.170 236.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1214.070 265.365 1217.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.070 10.640 1257.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1294.070 10.640 1297.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1334.070 10.640 1337.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.070 10.640 1377.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.070 10.640 1417.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.070 1046.620 1417.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.070 10.640 1457.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.070 1046.620 1457.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1494.070 10.640 1497.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1494.070 1046.620 1497.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.070 10.640 1537.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.070 1046.620 1537.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1574.070 10.640 1577.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1574.070 1046.620 1577.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.070 10.640 1617.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.070 1047.240 1617.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.070 10.640 1657.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.070 1047.240 1657.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1694.070 10.640 1697.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1694.070 1046.620 1697.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1734.070 10.640 1737.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1734.070 1046.620 1737.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.070 10.640 1777.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.070 1046.620 1777.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.070 10.640 1817.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.070 1047.240 1817.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1854.070 10.640 1857.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1854.070 1047.240 1857.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.070 10.640 1897.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.070 1046.620 1897.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.070 10.640 1937.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.070 1046.620 1937.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1974.070 10.640 1977.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1974.070 1046.620 1977.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2014.070 10.640 2017.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2014.070 1046.620 2017.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2054.070 10.640 2057.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2054.070 1047.240 2057.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.070 10.640 2097.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.070 10.640 2137.170 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.070 10.640 2177.170 1488.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.430 2194.440 22.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 59.430 2194.440 62.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 99.430 2194.440 102.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 139.430 2194.440 142.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.430 2194.440 182.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 219.430 2194.440 222.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 259.430 2194.440 262.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 299.430 2194.440 302.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 339.430 2194.440 342.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 379.430 2194.440 382.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 419.430 2194.440 422.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 459.430 2194.440 462.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 499.430 2194.440 502.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 539.430 2194.440 542.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 579.430 2194.440 582.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 619.430 2194.440 622.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 659.430 2194.440 662.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 699.430 2194.440 702.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 739.430 2194.440 742.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 779.430 2194.440 782.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 819.430 2194.440 822.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 859.430 2194.440 862.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 899.430 2194.440 902.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 939.430 2194.440 942.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 979.430 2194.440 982.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1019.430 2194.440 1022.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1059.430 2194.440 1062.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1099.430 2194.440 1102.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1139.430 2194.440 1142.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1179.430 2194.440 1182.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1219.430 2194.440 1222.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1259.430 2194.440 1262.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1299.430 2194.440 1302.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1339.430 2194.440 1342.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1379.430 2194.440 1382.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1419.430 2194.440 1422.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1459.430 2194.440 1462.530 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.970 10.640 52.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.970 10.640 92.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.970 1046.620 92.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.970 10.640 132.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.970 1046.620 132.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.970 10.640 172.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.970 1046.620 172.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 10.640 212.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 1046.620 212.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.970 10.640 252.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.970 1046.620 252.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 10.640 292.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 1046.960 292.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.970 10.640 332.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.970 1046.960 332.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1046.620 372.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 10.640 412.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 1046.620 412.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.970 10.640 452.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.970 1046.620 452.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.970 10.640 492.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.970 1046.620 492.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 528.970 10.640 532.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 528.970 1046.960 532.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 10.640 572.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 1046.620 572.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 10.640 612.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 1046.620 612.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.970 10.640 652.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.970 1046.620 652.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 688.970 10.640 692.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 688.970 1046.960 692.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 10.640 732.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1046.620 732.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 768.970 10.640 772.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 768.970 1046.620 772.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 10.640 812.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.970 10.640 852.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 888.970 10.640 892.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 928.970 10.640 932.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 968.970 10.640 972.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.970 10.640 1012.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1048.970 10.640 1052.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 10.640 1092.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.970 10.640 1132.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1168.970 10.640 1172.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.970 10.640 1212.070 189.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.970 273.940 1212.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1248.970 10.640 1252.070 189.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1248.970 273.940 1252.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1288.970 10.640 1292.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1328.970 10.640 1332.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1368.970 10.640 1372.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 10.640 1412.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 1046.620 1412.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 10.640 1452.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 1046.620 1452.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1488.970 10.640 1492.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1488.970 1046.620 1492.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1528.970 10.640 1532.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1528.970 1046.620 1532.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1568.970 10.640 1572.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1568.970 1046.620 1572.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.970 10.640 1612.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.970 1046.620 1612.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1648.970 10.640 1652.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1648.970 1046.620 1652.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 10.640 1692.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 1046.960 1692.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1728.970 10.640 1732.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1728.970 1046.960 1732.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.970 10.640 1772.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.970 1046.620 1772.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 10.640 1812.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 1046.620 1812.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1848.970 10.640 1852.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1848.970 1046.620 1852.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1888.970 10.640 1892.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1888.970 1046.960 1892.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1928.970 10.640 1932.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1928.970 1046.960 1932.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 10.640 1972.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 1046.620 1972.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.970 10.640 2012.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.970 1046.620 2012.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2048.970 10.640 2052.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2048.970 1046.620 2052.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2088.970 10.640 2092.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2088.970 1046.620 2092.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2128.970 10.640 2132.070 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 10.640 2172.070 1488.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 14.330 2194.440 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 54.330 2194.440 57.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 94.330 2194.440 97.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 134.330 2194.440 137.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 174.330 2194.440 177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 214.330 2194.440 217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 254.330 2194.440 257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 294.330 2194.440 297.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 334.330 2194.440 337.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 374.330 2194.440 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 414.330 2194.440 417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 454.330 2194.440 457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 494.330 2194.440 497.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 534.330 2194.440 537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 574.330 2194.440 577.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 614.330 2194.440 617.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 654.330 2194.440 657.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 694.330 2194.440 697.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 734.330 2194.440 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 774.330 2194.440 777.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 814.330 2194.440 817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 854.330 2194.440 857.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 894.330 2194.440 897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 934.330 2194.440 937.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 974.330 2194.440 977.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1014.330 2194.440 1017.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1054.330 2194.440 1057.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1094.330 2194.440 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1134.330 2194.440 1137.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1174.330 2194.440 1177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1214.330 2194.440 1217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1254.330 2194.440 1257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1294.330 2194.440 1297.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1334.330 2194.440 1337.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1374.330 2194.440 1377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1414.330 2194.440 1417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1454.330 2194.440 1457.430 ;
    END
  END VPWR
  PIN gpio_dm0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 43.560 2200.000 44.160 ;
    END
  END gpio_dm0[0]
  PIN gpio_dm0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1022.760 2200.000 1023.360 ;
    END
  END gpio_dm0[10]
  PIN gpio_dm0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1120.680 2200.000 1121.280 ;
    END
  END gpio_dm0[11]
  PIN gpio_dm0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1218.600 2200.000 1219.200 ;
    END
  END gpio_dm0[12]
  PIN gpio_dm0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1316.520 2200.000 1317.120 ;
    END
  END gpio_dm0[13]
  PIN gpio_dm0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1414.440 2200.000 1415.040 ;
    END
  END gpio_dm0[14]
  PIN gpio_dm0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2121.610 1497.600 2121.890 1500.000 ;
    END
  END gpio_dm0[15]
  PIN gpio_dm0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1878.730 1497.600 1879.010 1500.000 ;
    END
  END gpio_dm0[16]
  PIN gpio_dm0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1635.850 1497.600 1636.130 1500.000 ;
    END
  END gpio_dm0[17]
  PIN gpio_dm0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1392.970 1497.600 1393.250 1500.000 ;
    END
  END gpio_dm0[18]
  PIN gpio_dm0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1150.090 1497.600 1150.370 1500.000 ;
    END
  END gpio_dm0[19]
  PIN gpio_dm0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 141.480 2200.000 142.080 ;
    END
  END gpio_dm0[1]
  PIN gpio_dm0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 907.210 1497.600 907.490 1500.000 ;
    END
  END gpio_dm0[20]
  PIN gpio_dm0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 664.330 1497.600 664.610 1500.000 ;
    END
  END gpio_dm0[21]
  PIN gpio_dm0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 421.450 1497.600 421.730 1500.000 ;
    END
  END gpio_dm0[22]
  PIN gpio_dm0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 178.570 1497.600 178.850 1500.000 ;
    END
  END gpio_dm0[23]
  PIN gpio_dm0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1414.440 2.400 1415.040 ;
    END
  END gpio_dm0[24]
  PIN gpio_dm0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1316.520 2.400 1317.120 ;
    END
  END gpio_dm0[25]
  PIN gpio_dm0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1218.600 2.400 1219.200 ;
    END
  END gpio_dm0[26]
  PIN gpio_dm0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.680 2.400 1121.280 ;
    END
  END gpio_dm0[27]
  PIN gpio_dm0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.760 2.400 1023.360 ;
    END
  END gpio_dm0[28]
  PIN gpio_dm0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 2.400 925.440 ;
    END
  END gpio_dm0[29]
  PIN gpio_dm0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 239.400 2200.000 240.000 ;
    END
  END gpio_dm0[2]
  PIN gpio_dm0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.920 2.400 827.520 ;
    END
  END gpio_dm0[30]
  PIN gpio_dm0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 2.400 729.600 ;
    END
  END gpio_dm0[31]
  PIN gpio_dm0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 2.400 631.680 ;
    END
  END gpio_dm0[32]
  PIN gpio_dm0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 2.400 533.760 ;
    END
  END gpio_dm0[33]
  PIN gpio_dm0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 2.400 435.840 ;
    END
  END gpio_dm0[34]
  PIN gpio_dm0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 2.400 337.920 ;
    END
  END gpio_dm0[35]
  PIN gpio_dm0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 2.400 240.000 ;
    END
  END gpio_dm0[36]
  PIN gpio_dm0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 2.400 142.080 ;
    END
  END gpio_dm0[37]
  PIN gpio_dm0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 2.400 ;
    END
  END gpio_dm0[38]
  PIN gpio_dm0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 2.400 ;
    END
  END gpio_dm0[39]
  PIN gpio_dm0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 337.320 2200.000 337.920 ;
    END
  END gpio_dm0[3]
  PIN gpio_dm0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 2.400 ;
    END
  END gpio_dm0[40]
  PIN gpio_dm0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 2.400 ;
    END
  END gpio_dm0[41]
  PIN gpio_dm0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1099.490 0.000 1099.770 2.400 ;
    END
  END gpio_dm0[42]
  PIN gpio_dm0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1347.890 0.000 1348.170 2.400 ;
    END
  END gpio_dm0[43]
  PIN gpio_dm0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 435.240 2200.000 435.840 ;
    END
  END gpio_dm0[4]
  PIN gpio_dm0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 533.160 2200.000 533.760 ;
    END
  END gpio_dm0[5]
  PIN gpio_dm0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 631.080 2200.000 631.680 ;
    END
  END gpio_dm0[6]
  PIN gpio_dm0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 729.000 2200.000 729.600 ;
    END
  END gpio_dm0[7]
  PIN gpio_dm0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 826.920 2200.000 827.520 ;
    END
  END gpio_dm0[8]
  PIN gpio_dm0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 924.840 2200.000 925.440 ;
    END
  END gpio_dm0[9]
  PIN gpio_dm1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 35.400 2200.000 36.000 ;
    END
  END gpio_dm1[0]
  PIN gpio_dm1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1014.600 2200.000 1015.200 ;
    END
  END gpio_dm1[10]
  PIN gpio_dm1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1112.520 2200.000 1113.120 ;
    END
  END gpio_dm1[11]
  PIN gpio_dm1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1210.440 2200.000 1211.040 ;
    END
  END gpio_dm1[12]
  PIN gpio_dm1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1308.360 2200.000 1308.960 ;
    END
  END gpio_dm1[13]
  PIN gpio_dm1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1406.280 2200.000 1406.880 ;
    END
  END gpio_dm1[14]
  PIN gpio_dm1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2141.850 1497.600 2142.130 1500.000 ;
    END
  END gpio_dm1[15]
  PIN gpio_dm1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1898.970 1497.600 1899.250 1500.000 ;
    END
  END gpio_dm1[16]
  PIN gpio_dm1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1656.090 1497.600 1656.370 1500.000 ;
    END
  END gpio_dm1[17]
  PIN gpio_dm1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1413.210 1497.600 1413.490 1500.000 ;
    END
  END gpio_dm1[18]
  PIN gpio_dm1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1170.330 1497.600 1170.610 1500.000 ;
    END
  END gpio_dm1[19]
  PIN gpio_dm1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 133.320 2200.000 133.920 ;
    END
  END gpio_dm1[1]
  PIN gpio_dm1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 927.450 1497.600 927.730 1500.000 ;
    END
  END gpio_dm1[20]
  PIN gpio_dm1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 684.570 1497.600 684.850 1500.000 ;
    END
  END gpio_dm1[21]
  PIN gpio_dm1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 441.690 1497.600 441.970 1500.000 ;
    END
  END gpio_dm1[22]
  PIN gpio_dm1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 198.810 1497.600 199.090 1500.000 ;
    END
  END gpio_dm1[23]
  PIN gpio_dm1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1422.600 2.400 1423.200 ;
    END
  END gpio_dm1[24]
  PIN gpio_dm1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.680 2.400 1325.280 ;
    END
  END gpio_dm1[25]
  PIN gpio_dm1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1226.760 2.400 1227.360 ;
    END
  END gpio_dm1[26]
  PIN gpio_dm1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 2.400 1129.440 ;
    END
  END gpio_dm1[27]
  PIN gpio_dm1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.920 2.400 1031.520 ;
    END
  END gpio_dm1[28]
  PIN gpio_dm1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 2.400 933.600 ;
    END
  END gpio_dm1[29]
  PIN gpio_dm1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 231.240 2200.000 231.840 ;
    END
  END gpio_dm1[2]
  PIN gpio_dm1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 2.400 835.680 ;
    END
  END gpio_dm1[30]
  PIN gpio_dm1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 2.400 737.760 ;
    END
  END gpio_dm1[31]
  PIN gpio_dm1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 2.400 639.840 ;
    END
  END gpio_dm1[32]
  PIN gpio_dm1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 2.400 541.920 ;
    END
  END gpio_dm1[33]
  PIN gpio_dm1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 2.400 444.000 ;
    END
  END gpio_dm1[34]
  PIN gpio_dm1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 2.400 346.080 ;
    END
  END gpio_dm1[35]
  PIN gpio_dm1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 2.400 248.160 ;
    END
  END gpio_dm1[36]
  PIN gpio_dm1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 2.400 150.240 ;
    END
  END gpio_dm1[37]
  PIN gpio_dm1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 2.400 ;
    END
  END gpio_dm1[38]
  PIN gpio_dm1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 2.400 ;
    END
  END gpio_dm1[39]
  PIN gpio_dm1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 329.160 2200.000 329.760 ;
    END
  END gpio_dm1[3]
  PIN gpio_dm1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 2.400 ;
    END
  END gpio_dm1[40]
  PIN gpio_dm1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 2.400 ;
    END
  END gpio_dm1[41]
  PIN gpio_dm1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 2.400 ;
    END
  END gpio_dm1[42]
  PIN gpio_dm1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1327.190 0.000 1327.470 2.400 ;
    END
  END gpio_dm1[43]
  PIN gpio_dm1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 427.080 2200.000 427.680 ;
    END
  END gpio_dm1[4]
  PIN gpio_dm1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 525.000 2200.000 525.600 ;
    END
  END gpio_dm1[5]
  PIN gpio_dm1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 622.920 2200.000 623.520 ;
    END
  END gpio_dm1[6]
  PIN gpio_dm1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 720.840 2200.000 721.440 ;
    END
  END gpio_dm1[7]
  PIN gpio_dm1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 818.760 2200.000 819.360 ;
    END
  END gpio_dm1[8]
  PIN gpio_dm1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 916.680 2200.000 917.280 ;
    END
  END gpio_dm1[9]
  PIN gpio_dm2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 59.880 2200.000 60.480 ;
    END
  END gpio_dm2[0]
  PIN gpio_dm2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1039.080 2200.000 1039.680 ;
    END
  END gpio_dm2[10]
  PIN gpio_dm2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1137.000 2200.000 1137.600 ;
    END
  END gpio_dm2[11]
  PIN gpio_dm2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1234.920 2200.000 1235.520 ;
    END
  END gpio_dm2[12]
  PIN gpio_dm2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1332.840 2200.000 1333.440 ;
    END
  END gpio_dm2[13]
  PIN gpio_dm2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1430.760 2200.000 1431.360 ;
    END
  END gpio_dm2[14]
  PIN gpio_dm2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2081.130 1497.600 2081.410 1500.000 ;
    END
  END gpio_dm2[15]
  PIN gpio_dm2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1838.250 1497.600 1838.530 1500.000 ;
    END
  END gpio_dm2[16]
  PIN gpio_dm2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1595.370 1497.600 1595.650 1500.000 ;
    END
  END gpio_dm2[17]
  PIN gpio_dm2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1352.490 1497.600 1352.770 1500.000 ;
    END
  END gpio_dm2[18]
  PIN gpio_dm2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1109.610 1497.600 1109.890 1500.000 ;
    END
  END gpio_dm2[19]
  PIN gpio_dm2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 157.800 2200.000 158.400 ;
    END
  END gpio_dm2[1]
  PIN gpio_dm2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 866.730 1497.600 867.010 1500.000 ;
    END
  END gpio_dm2[20]
  PIN gpio_dm2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 623.850 1497.600 624.130 1500.000 ;
    END
  END gpio_dm2[21]
  PIN gpio_dm2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 380.970 1497.600 381.250 1500.000 ;
    END
  END gpio_dm2[22]
  PIN gpio_dm2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 138.090 1497.600 138.370 1500.000 ;
    END
  END gpio_dm2[23]
  PIN gpio_dm2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1398.120 2.400 1398.720 ;
    END
  END gpio_dm2[24]
  PIN gpio_dm2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.200 2.400 1300.800 ;
    END
  END gpio_dm2[25]
  PIN gpio_dm2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.280 2.400 1202.880 ;
    END
  END gpio_dm2[26]
  PIN gpio_dm2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1104.360 2.400 1104.960 ;
    END
  END gpio_dm2[27]
  PIN gpio_dm2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 2.400 1007.040 ;
    END
  END gpio_dm2[28]
  PIN gpio_dm2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 2.400 909.120 ;
    END
  END gpio_dm2[29]
  PIN gpio_dm2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 255.720 2200.000 256.320 ;
    END
  END gpio_dm2[2]
  PIN gpio_dm2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 2.400 811.200 ;
    END
  END gpio_dm2[30]
  PIN gpio_dm2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 2.400 713.280 ;
    END
  END gpio_dm2[31]
  PIN gpio_dm2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 2.400 615.360 ;
    END
  END gpio_dm2[32]
  PIN gpio_dm2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 2.400 517.440 ;
    END
  END gpio_dm2[33]
  PIN gpio_dm2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 2.400 419.520 ;
    END
  END gpio_dm2[34]
  PIN gpio_dm2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 2.400 321.600 ;
    END
  END gpio_dm2[35]
  PIN gpio_dm2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 2.400 223.680 ;
    END
  END gpio_dm2[36]
  PIN gpio_dm2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 2.400 125.760 ;
    END
  END gpio_dm2[37]
  PIN gpio_dm2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 2.400 ;
    END
  END gpio_dm2[38]
  PIN gpio_dm2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 2.400 ;
    END
  END gpio_dm2[39]
  PIN gpio_dm2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 353.640 2200.000 354.240 ;
    END
  END gpio_dm2[3]
  PIN gpio_dm2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 2.400 ;
    END
  END gpio_dm2[40]
  PIN gpio_dm2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 2.400 ;
    END
  END gpio_dm2[41]
  PIN gpio_dm2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1140.890 0.000 1141.170 2.400 ;
    END
  END gpio_dm2[42]
  PIN gpio_dm2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1389.290 0.000 1389.570 2.400 ;
    END
  END gpio_dm2[43]
  PIN gpio_dm2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 451.560 2200.000 452.160 ;
    END
  END gpio_dm2[4]
  PIN gpio_dm2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 549.480 2200.000 550.080 ;
    END
  END gpio_dm2[5]
  PIN gpio_dm2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 647.400 2200.000 648.000 ;
    END
  END gpio_dm2[6]
  PIN gpio_dm2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 745.320 2200.000 745.920 ;
    END
  END gpio_dm2[7]
  PIN gpio_dm2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 843.240 2200.000 843.840 ;
    END
  END gpio_dm2[8]
  PIN gpio_dm2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 941.160 2200.000 941.760 ;
    END
  END gpio_dm2[9]
  PIN gpio_ib_mode_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 84.360 2200.000 84.960 ;
    END
  END gpio_ib_mode_sel[0]
  PIN gpio_ib_mode_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1063.560 2200.000 1064.160 ;
    END
  END gpio_ib_mode_sel[10]
  PIN gpio_ib_mode_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1161.480 2200.000 1162.080 ;
    END
  END gpio_ib_mode_sel[11]
  PIN gpio_ib_mode_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1259.400 2200.000 1260.000 ;
    END
  END gpio_ib_mode_sel[12]
  PIN gpio_ib_mode_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1357.320 2200.000 1357.920 ;
    END
  END gpio_ib_mode_sel[13]
  PIN gpio_ib_mode_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1455.240 2200.000 1455.840 ;
    END
  END gpio_ib_mode_sel[14]
  PIN gpio_ib_mode_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2020.410 1497.600 2020.690 1500.000 ;
    END
  END gpio_ib_mode_sel[15]
  PIN gpio_ib_mode_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1777.530 1497.600 1777.810 1500.000 ;
    END
  END gpio_ib_mode_sel[16]
  PIN gpio_ib_mode_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1534.650 1497.600 1534.930 1500.000 ;
    END
  END gpio_ib_mode_sel[17]
  PIN gpio_ib_mode_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1291.770 1497.600 1292.050 1500.000 ;
    END
  END gpio_ib_mode_sel[18]
  PIN gpio_ib_mode_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1048.890 1497.600 1049.170 1500.000 ;
    END
  END gpio_ib_mode_sel[19]
  PIN gpio_ib_mode_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 182.280 2200.000 182.880 ;
    END
  END gpio_ib_mode_sel[1]
  PIN gpio_ib_mode_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 806.010 1497.600 806.290 1500.000 ;
    END
  END gpio_ib_mode_sel[20]
  PIN gpio_ib_mode_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 563.130 1497.600 563.410 1500.000 ;
    END
  END gpio_ib_mode_sel[21]
  PIN gpio_ib_mode_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 320.250 1497.600 320.530 1500.000 ;
    END
  END gpio_ib_mode_sel[22]
  PIN gpio_ib_mode_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 77.370 1497.600 77.650 1500.000 ;
    END
  END gpio_ib_mode_sel[23]
  PIN gpio_ib_mode_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 2.400 1374.240 ;
    END
  END gpio_ib_mode_sel[24]
  PIN gpio_ib_mode_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.720 2.400 1276.320 ;
    END
  END gpio_ib_mode_sel[25]
  PIN gpio_ib_mode_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.800 2.400 1178.400 ;
    END
  END gpio_ib_mode_sel[26]
  PIN gpio_ib_mode_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1079.880 2.400 1080.480 ;
    END
  END gpio_ib_mode_sel[27]
  PIN gpio_ib_mode_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.960 2.400 982.560 ;
    END
  END gpio_ib_mode_sel[28]
  PIN gpio_ib_mode_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 2.400 884.640 ;
    END
  END gpio_ib_mode_sel[29]
  PIN gpio_ib_mode_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 280.200 2200.000 280.800 ;
    END
  END gpio_ib_mode_sel[2]
  PIN gpio_ib_mode_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 2.400 786.720 ;
    END
  END gpio_ib_mode_sel[30]
  PIN gpio_ib_mode_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 2.400 688.800 ;
    END
  END gpio_ib_mode_sel[31]
  PIN gpio_ib_mode_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 2.400 590.880 ;
    END
  END gpio_ib_mode_sel[32]
  PIN gpio_ib_mode_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 2.400 492.960 ;
    END
  END gpio_ib_mode_sel[33]
  PIN gpio_ib_mode_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 2.400 395.040 ;
    END
  END gpio_ib_mode_sel[34]
  PIN gpio_ib_mode_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 2.400 297.120 ;
    END
  END gpio_ib_mode_sel[35]
  PIN gpio_ib_mode_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 2.400 199.200 ;
    END
  END gpio_ib_mode_sel[36]
  PIN gpio_ib_mode_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END gpio_ib_mode_sel[37]
  PIN gpio_ib_mode_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 2.400 ;
    END
  END gpio_ib_mode_sel[38]
  PIN gpio_ib_mode_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 2.400 ;
    END
  END gpio_ib_mode_sel[39]
  PIN gpio_ib_mode_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 378.120 2200.000 378.720 ;
    END
  END gpio_ib_mode_sel[3]
  PIN gpio_ib_mode_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 2.400 ;
    END
  END gpio_ib_mode_sel[40]
  PIN gpio_ib_mode_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 954.590 0.000 954.870 2.400 ;
    END
  END gpio_ib_mode_sel[41]
  PIN gpio_ib_mode_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1202.990 0.000 1203.270 2.400 ;
    END
  END gpio_ib_mode_sel[42]
  PIN gpio_ib_mode_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1451.390 0.000 1451.670 2.400 ;
    END
  END gpio_ib_mode_sel[43]
  PIN gpio_ib_mode_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 476.040 2200.000 476.640 ;
    END
  END gpio_ib_mode_sel[4]
  PIN gpio_ib_mode_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 573.960 2200.000 574.560 ;
    END
  END gpio_ib_mode_sel[5]
  PIN gpio_ib_mode_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 671.880 2200.000 672.480 ;
    END
  END gpio_ib_mode_sel[6]
  PIN gpio_ib_mode_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 769.800 2200.000 770.400 ;
    END
  END gpio_ib_mode_sel[7]
  PIN gpio_ib_mode_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 867.720 2200.000 868.320 ;
    END
  END gpio_ib_mode_sel[8]
  PIN gpio_ib_mode_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 965.640 2200.000 966.240 ;
    END
  END gpio_ib_mode_sel[9]
  PIN gpio_ieb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 51.720 2200.000 52.320 ;
    END
  END gpio_ieb[0]
  PIN gpio_ieb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1030.920 2200.000 1031.520 ;
    END
  END gpio_ieb[10]
  PIN gpio_ieb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1128.840 2200.000 1129.440 ;
    END
  END gpio_ieb[11]
  PIN gpio_ieb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1226.760 2200.000 1227.360 ;
    END
  END gpio_ieb[12]
  PIN gpio_ieb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1324.680 2200.000 1325.280 ;
    END
  END gpio_ieb[13]
  PIN gpio_ieb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1422.600 2200.000 1423.200 ;
    END
  END gpio_ieb[14]
  PIN gpio_ieb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2101.370 1497.600 2101.650 1500.000 ;
    END
  END gpio_ieb[15]
  PIN gpio_ieb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1858.490 1497.600 1858.770 1500.000 ;
    END
  END gpio_ieb[16]
  PIN gpio_ieb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1615.610 1497.600 1615.890 1500.000 ;
    END
  END gpio_ieb[17]
  PIN gpio_ieb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1372.730 1497.600 1373.010 1500.000 ;
    END
  END gpio_ieb[18]
  PIN gpio_ieb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1129.850 1497.600 1130.130 1500.000 ;
    END
  END gpio_ieb[19]
  PIN gpio_ieb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 149.640 2200.000 150.240 ;
    END
  END gpio_ieb[1]
  PIN gpio_ieb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 886.970 1497.600 887.250 1500.000 ;
    END
  END gpio_ieb[20]
  PIN gpio_ieb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 644.090 1497.600 644.370 1500.000 ;
    END
  END gpio_ieb[21]
  PIN gpio_ieb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 401.210 1497.600 401.490 1500.000 ;
    END
  END gpio_ieb[22]
  PIN gpio_ieb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 158.330 1497.600 158.610 1500.000 ;
    END
  END gpio_ieb[23]
  PIN gpio_ieb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1406.280 2.400 1406.880 ;
    END
  END gpio_ieb[24]
  PIN gpio_ieb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1308.360 2.400 1308.960 ;
    END
  END gpio_ieb[25]
  PIN gpio_ieb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1210.440 2.400 1211.040 ;
    END
  END gpio_ieb[26]
  PIN gpio_ieb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1112.520 2.400 1113.120 ;
    END
  END gpio_ieb[27]
  PIN gpio_ieb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1014.600 2.400 1015.200 ;
    END
  END gpio_ieb[28]
  PIN gpio_ieb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 2.400 917.280 ;
    END
  END gpio_ieb[29]
  PIN gpio_ieb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 247.560 2200.000 248.160 ;
    END
  END gpio_ieb[2]
  PIN gpio_ieb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 2.400 819.360 ;
    END
  END gpio_ieb[30]
  PIN gpio_ieb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 2.400 721.440 ;
    END
  END gpio_ieb[31]
  PIN gpio_ieb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 2.400 623.520 ;
    END
  END gpio_ieb[32]
  PIN gpio_ieb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 2.400 525.600 ;
    END
  END gpio_ieb[33]
  PIN gpio_ieb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 2.400 427.680 ;
    END
  END gpio_ieb[34]
  PIN gpio_ieb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 2.400 329.760 ;
    END
  END gpio_ieb[35]
  PIN gpio_ieb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 2.400 231.840 ;
    END
  END gpio_ieb[36]
  PIN gpio_ieb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 2.400 133.920 ;
    END
  END gpio_ieb[37]
  PIN gpio_ieb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 2.400 ;
    END
  END gpio_ieb[38]
  PIN gpio_ieb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 2.400 ;
    END
  END gpio_ieb[39]
  PIN gpio_ieb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 345.480 2200.000 346.080 ;
    END
  END gpio_ieb[3]
  PIN gpio_ieb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 2.400 ;
    END
  END gpio_ieb[40]
  PIN gpio_ieb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 2.400 ;
    END
  END gpio_ieb[41]
  PIN gpio_ieb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 2.400 ;
    END
  END gpio_ieb[42]
  PIN gpio_ieb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 2.400 ;
    END
  END gpio_ieb[43]
  PIN gpio_ieb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 443.400 2200.000 444.000 ;
    END
  END gpio_ieb[4]
  PIN gpio_ieb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 541.320 2200.000 541.920 ;
    END
  END gpio_ieb[5]
  PIN gpio_ieb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 639.240 2200.000 639.840 ;
    END
  END gpio_ieb[6]
  PIN gpio_ieb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 737.160 2200.000 737.760 ;
    END
  END gpio_ieb[7]
  PIN gpio_ieb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 835.080 2200.000 835.680 ;
    END
  END gpio_ieb[8]
  PIN gpio_ieb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 933.000 2200.000 933.600 ;
    END
  END gpio_ieb[9]
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 19.080 2200.000 19.680 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 998.280 2200.000 998.880 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1096.200 2200.000 1096.800 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1194.120 2200.000 1194.720 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1292.040 2200.000 1292.640 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1389.960 2200.000 1390.560 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2182.330 1497.600 2182.610 1500.000 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1939.450 1497.600 1939.730 1500.000 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1696.570 1497.600 1696.850 1500.000 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1453.690 1497.600 1453.970 1500.000 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1210.810 1497.600 1211.090 1500.000 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 117.000 2200.000 117.600 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 967.930 1497.600 968.210 1500.000 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 725.050 1497.600 725.330 1500.000 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 482.170 1497.600 482.450 1500.000 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 239.290 1497.600 239.570 1500.000 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.920 2.400 1439.520 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1341.000 2.400 1341.600 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 2.400 1243.680 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 2.400 1145.760 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 2.400 1047.840 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 949.320 2.400 949.920 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 214.920 2200.000 215.520 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 2.400 852.000 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 753.480 2.400 754.080 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 2.400 656.160 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 2.400 558.240 ;
    END
  END gpio_in[33]
  PIN gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 2.400 460.320 ;
    END
  END gpio_in[34]
  PIN gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 2.400 362.400 ;
    END
  END gpio_in[35]
  PIN gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 2.400 264.480 ;
    END
  END gpio_in[36]
  PIN gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 2.400 166.560 ;
    END
  END gpio_in[37]
  PIN gpio_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.400 ;
    END
  END gpio_in[38]
  PIN gpio_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 2.400 ;
    END
  END gpio_in[39]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 312.840 2200.000 313.440 ;
    END
  END gpio_in[3]
  PIN gpio_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 2.400 ;
    END
  END gpio_in[40]
  PIN gpio_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 2.400 ;
    END
  END gpio_in[41]
  PIN gpio_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 2.400 ;
    END
  END gpio_in[42]
  PIN gpio_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1285.790 0.000 1286.070 2.400 ;
    END
  END gpio_in[43]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 410.760 2200.000 411.360 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 508.680 2200.000 509.280 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 606.600 2200.000 607.200 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 704.520 2200.000 705.120 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 802.440 2200.000 803.040 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 900.360 2200.000 900.960 ;
    END
  END gpio_in[9]
  PIN gpio_loopback_one[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2197.600 100.680 2200.000 101.280 ;
    END
  END gpio_loopback_one[0]
  PIN gpio_loopback_one[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1079.880 2200.000 1080.480 ;
    END
  END gpio_loopback_one[10]
  PIN gpio_loopback_one[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1177.800 2200.000 1178.400 ;
    END
  END gpio_loopback_one[11]
  PIN gpio_loopback_one[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1275.720 2200.000 1276.320 ;
    END
  END gpio_loopback_one[12]
  PIN gpio_loopback_one[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1373.640 2200.000 1374.240 ;
    END
  END gpio_loopback_one[13]
  PIN gpio_loopback_one[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1471.560 2200.000 1472.160 ;
    END
  END gpio_loopback_one[14]
  PIN gpio_loopback_one[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1979.930 1497.600 1980.210 1500.000 ;
    END
  END gpio_loopback_one[15]
  PIN gpio_loopback_one[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.050 1497.600 1737.330 1500.000 ;
    END
  END gpio_loopback_one[16]
  PIN gpio_loopback_one[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 1497.600 1494.450 1500.000 ;
    END
  END gpio_loopback_one[17]
  PIN gpio_loopback_one[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.290 1497.600 1251.570 1500.000 ;
    END
  END gpio_loopback_one[18]
  PIN gpio_loopback_one[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 1497.600 1008.690 1500.000 ;
    END
  END gpio_loopback_one[19]
  PIN gpio_loopback_one[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 198.600 2200.000 199.200 ;
    END
  END gpio_loopback_one[1]
  PIN gpio_loopback_one[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 1497.600 765.810 1500.000 ;
    END
  END gpio_loopback_one[20]
  PIN gpio_loopback_one[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 1497.600 522.930 1500.000 ;
    END
  END gpio_loopback_one[21]
  PIN gpio_loopback_one[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 1497.600 280.050 1500.000 ;
    END
  END gpio_loopback_one[22]
  PIN gpio_loopback_one[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 1497.600 37.170 1500.000 ;
    END
  END gpio_loopback_one[23]
  PIN gpio_loopback_one[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1357.320 2.400 1357.920 ;
    END
  END gpio_loopback_one[24]
  PIN gpio_loopback_one[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1259.400 2.400 1260.000 ;
    END
  END gpio_loopback_one[25]
  PIN gpio_loopback_one[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1161.480 2.400 1162.080 ;
    END
  END gpio_loopback_one[26]
  PIN gpio_loopback_one[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1063.560 2.400 1064.160 ;
    END
  END gpio_loopback_one[27]
  PIN gpio_loopback_one[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 2.400 966.240 ;
    END
  END gpio_loopback_one[28]
  PIN gpio_loopback_one[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 2.400 868.320 ;
    END
  END gpio_loopback_one[29]
  PIN gpio_loopback_one[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 296.520 2200.000 297.120 ;
    END
  END gpio_loopback_one[2]
  PIN gpio_loopback_one[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 2.400 770.400 ;
    END
  END gpio_loopback_one[30]
  PIN gpio_loopback_one[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 2.400 672.480 ;
    END
  END gpio_loopback_one[31]
  PIN gpio_loopback_one[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 2.400 574.560 ;
    END
  END gpio_loopback_one[32]
  PIN gpio_loopback_one[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 2.400 476.640 ;
    END
  END gpio_loopback_one[33]
  PIN gpio_loopback_one[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 2.400 378.720 ;
    END
  END gpio_loopback_one[34]
  PIN gpio_loopback_one[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 2.400 280.800 ;
    END
  END gpio_loopback_one[35]
  PIN gpio_loopback_one[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 2.400 182.880 ;
    END
  END gpio_loopback_one[36]
  PIN gpio_loopback_one[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 2.400 84.960 ;
    END
  END gpio_loopback_one[37]
  PIN gpio_loopback_one[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 2.400 ;
    END
  END gpio_loopback_one[38]
  PIN gpio_loopback_one[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 2.400 ;
    END
  END gpio_loopback_one[39]
  PIN gpio_loopback_one[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 394.440 2200.000 395.040 ;
    END
  END gpio_loopback_one[3]
  PIN gpio_loopback_one[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 2.400 ;
    END
  END gpio_loopback_one[40]
  PIN gpio_loopback_one[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 2.400 ;
    END
  END gpio_loopback_one[41]
  PIN gpio_loopback_one[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 0.000 1244.670 2.400 ;
    END
  END gpio_loopback_one[42]
  PIN gpio_loopback_one[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 0.000 1493.070 2.400 ;
    END
  END gpio_loopback_one[43]
  PIN gpio_loopback_one[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 492.360 2200.000 492.960 ;
    END
  END gpio_loopback_one[4]
  PIN gpio_loopback_one[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 590.280 2200.000 590.880 ;
    END
  END gpio_loopback_one[5]
  PIN gpio_loopback_one[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 688.200 2200.000 688.800 ;
    END
  END gpio_loopback_one[6]
  PIN gpio_loopback_one[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 786.120 2200.000 786.720 ;
    END
  END gpio_loopback_one[7]
  PIN gpio_loopback_one[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 884.040 2200.000 884.640 ;
    END
  END gpio_loopback_one[8]
  PIN gpio_loopback_one[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 981.960 2200.000 982.560 ;
    END
  END gpio_loopback_one[9]
  PIN gpio_loopback_zero[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2197.600 108.840 2200.000 109.440 ;
    END
  END gpio_loopback_zero[0]
  PIN gpio_loopback_zero[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1088.040 2200.000 1088.640 ;
    END
  END gpio_loopback_zero[10]
  PIN gpio_loopback_zero[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1185.960 2200.000 1186.560 ;
    END
  END gpio_loopback_zero[11]
  PIN gpio_loopback_zero[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1283.880 2200.000 1284.480 ;
    END
  END gpio_loopback_zero[12]
  PIN gpio_loopback_zero[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1381.800 2200.000 1382.400 ;
    END
  END gpio_loopback_zero[13]
  PIN gpio_loopback_zero[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1479.720 2200.000 1480.320 ;
    END
  END gpio_loopback_zero[14]
  PIN gpio_loopback_zero[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1959.690 1497.600 1959.970 1500.000 ;
    END
  END gpio_loopback_zero[15]
  PIN gpio_loopback_zero[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 1497.600 1717.090 1500.000 ;
    END
  END gpio_loopback_zero[16]
  PIN gpio_loopback_zero[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 1497.600 1474.210 1500.000 ;
    END
  END gpio_loopback_zero[17]
  PIN gpio_loopback_zero[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 1497.600 1231.330 1500.000 ;
    END
  END gpio_loopback_zero[18]
  PIN gpio_loopback_zero[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 1497.600 988.450 1500.000 ;
    END
  END gpio_loopback_zero[19]
  PIN gpio_loopback_zero[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2197.600 206.760 2200.000 207.360 ;
    END
  END gpio_loopback_zero[1]
  PIN gpio_loopback_zero[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 1497.600 745.570 1500.000 ;
    END
  END gpio_loopback_zero[20]
  PIN gpio_loopback_zero[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1497.600 502.690 1500.000 ;
    END
  END gpio_loopback_zero[21]
  PIN gpio_loopback_zero[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 1497.600 259.810 1500.000 ;
    END
  END gpio_loopback_zero[22]
  PIN gpio_loopback_zero[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 1497.600 16.930 1500.000 ;
    END
  END gpio_loopback_zero[23]
  PIN gpio_loopback_zero[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.160 2.400 1349.760 ;
    END
  END gpio_loopback_zero[24]
  PIN gpio_loopback_zero[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.240 2.400 1251.840 ;
    END
  END gpio_loopback_zero[25]
  PIN gpio_loopback_zero[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1153.320 2.400 1153.920 ;
    END
  END gpio_loopback_zero[26]
  PIN gpio_loopback_zero[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1055.400 2.400 1056.000 ;
    END
  END gpio_loopback_zero[27]
  PIN gpio_loopback_zero[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 957.480 2.400 958.080 ;
    END
  END gpio_loopback_zero[28]
  PIN gpio_loopback_zero[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 2.400 860.160 ;
    END
  END gpio_loopback_zero[29]
  PIN gpio_loopback_zero[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 304.680 2200.000 305.280 ;
    END
  END gpio_loopback_zero[2]
  PIN gpio_loopback_zero[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 2.400 762.240 ;
    END
  END gpio_loopback_zero[30]
  PIN gpio_loopback_zero[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 2.400 664.320 ;
    END
  END gpio_loopback_zero[31]
  PIN gpio_loopback_zero[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 2.400 566.400 ;
    END
  END gpio_loopback_zero[32]
  PIN gpio_loopback_zero[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 2.400 468.480 ;
    END
  END gpio_loopback_zero[33]
  PIN gpio_loopback_zero[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 2.400 370.560 ;
    END
  END gpio_loopback_zero[34]
  PIN gpio_loopback_zero[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 2.400 272.640 ;
    END
  END gpio_loopback_zero[35]
  PIN gpio_loopback_zero[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 2.400 174.720 ;
    END
  END gpio_loopback_zero[36]
  PIN gpio_loopback_zero[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 2.400 76.800 ;
    END
  END gpio_loopback_zero[37]
  PIN gpio_loopback_zero[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 2.400 ;
    END
  END gpio_loopback_zero[38]
  PIN gpio_loopback_zero[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 2.400 ;
    END
  END gpio_loopback_zero[39]
  PIN gpio_loopback_zero[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 402.600 2200.000 403.200 ;
    END
  END gpio_loopback_zero[3]
  PIN gpio_loopback_zero[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 2.400 ;
    END
  END gpio_loopback_zero[40]
  PIN gpio_loopback_zero[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 2.400 ;
    END
  END gpio_loopback_zero[41]
  PIN gpio_loopback_zero[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.090 0.000 1265.370 2.400 ;
    END
  END gpio_loopback_zero[42]
  PIN gpio_loopback_zero[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 0.000 1513.770 2.400 ;
    END
  END gpio_loopback_zero[43]
  PIN gpio_loopback_zero[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 500.520 2200.000 501.120 ;
    END
  END gpio_loopback_zero[4]
  PIN gpio_loopback_zero[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 598.440 2200.000 599.040 ;
    END
  END gpio_loopback_zero[5]
  PIN gpio_loopback_zero[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 696.360 2200.000 696.960 ;
    END
  END gpio_loopback_zero[6]
  PIN gpio_loopback_zero[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 794.280 2200.000 794.880 ;
    END
  END gpio_loopback_zero[7]
  PIN gpio_loopback_zero[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 892.200 2200.000 892.800 ;
    END
  END gpio_loopback_zero[8]
  PIN gpio_loopback_zero[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 990.120 2200.000 990.720 ;
    END
  END gpio_loopback_zero[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 92.520 2200.000 93.120 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1071.720 2200.000 1072.320 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1169.640 2200.000 1170.240 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1267.560 2200.000 1268.160 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1365.480 2200.000 1366.080 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1463.400 2200.000 1464.000 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2000.170 1497.600 2000.450 1500.000 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1757.290 1497.600 1757.570 1500.000 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1514.410 1497.600 1514.690 1500.000 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1271.530 1497.600 1271.810 1500.000 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1028.650 1497.600 1028.930 1500.000 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 190.440 2200.000 191.040 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 785.770 1497.600 786.050 1500.000 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 542.890 1497.600 543.170 1500.000 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 300.010 1497.600 300.290 1500.000 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 57.130 1497.600 57.410 1500.000 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1365.480 2.400 1366.080 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1267.560 2.400 1268.160 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 2.400 1170.240 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.720 2.400 1072.320 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.800 2.400 974.400 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 2.400 876.480 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 288.360 2200.000 288.960 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.960 2.400 778.560 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 2.400 680.640 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 2.400 582.720 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 2.400 484.800 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 2.400 386.880 ;
    END
  END gpio_oeb[34]
  PIN gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 2.400 288.960 ;
    END
  END gpio_oeb[35]
  PIN gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 2.400 191.040 ;
    END
  END gpio_oeb[36]
  PIN gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END gpio_oeb[37]
  PIN gpio_oeb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 2.400 ;
    END
  END gpio_oeb[38]
  PIN gpio_oeb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 2.400 ;
    END
  END gpio_oeb[39]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 386.280 2200.000 386.880 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 2.400 ;
    END
  END gpio_oeb[40]
  PIN gpio_oeb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 975.290 0.000 975.570 2.400 ;
    END
  END gpio_oeb[41]
  PIN gpio_oeb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 2.400 ;
    END
  END gpio_oeb[42]
  PIN gpio_oeb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1472.090 0.000 1472.370 2.400 ;
    END
  END gpio_oeb[43]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 484.200 2200.000 484.800 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 582.120 2200.000 582.720 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 680.040 2200.000 680.640 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 777.960 2200.000 778.560 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 875.880 2200.000 876.480 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 973.800 2200.000 974.400 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 68.040 2200.000 68.640 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1047.240 2200.000 1047.840 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1145.160 2200.000 1145.760 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1243.080 2200.000 1243.680 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1341.000 2200.000 1341.600 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1438.920 2200.000 1439.520 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2060.890 1497.600 2061.170 1500.000 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1818.010 1497.600 1818.290 1500.000 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1575.130 1497.600 1575.410 1500.000 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1332.250 1497.600 1332.530 1500.000 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1089.370 1497.600 1089.650 1500.000 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 165.960 2200.000 166.560 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 846.490 1497.600 846.770 1500.000 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 603.610 1497.600 603.890 1500.000 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 360.730 1497.600 361.010 1500.000 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 117.850 1497.600 118.130 1500.000 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1389.960 2.400 1390.560 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1292.040 2.400 1292.640 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 2.400 1194.720 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.200 2.400 1096.800 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 998.280 2.400 998.880 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 900.360 2.400 900.960 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 263.880 2200.000 264.480 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 2.400 803.040 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 2.400 705.120 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 2.400 607.200 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 2.400 509.280 ;
    END
  END gpio_out[33]
  PIN gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 2.400 411.360 ;
    END
  END gpio_out[34]
  PIN gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 2.400 313.440 ;
    END
  END gpio_out[35]
  PIN gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 2.400 215.520 ;
    END
  END gpio_out[36]
  PIN gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 2.400 117.600 ;
    END
  END gpio_out[37]
  PIN gpio_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 2.400 ;
    END
  END gpio_out[38]
  PIN gpio_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 2.400 ;
    END
  END gpio_out[39]
  PIN gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 361.800 2200.000 362.400 ;
    END
  END gpio_out[3]
  PIN gpio_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 664.790 0.000 665.070 2.400 ;
    END
  END gpio_out[40]
  PIN gpio_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 2.400 ;
    END
  END gpio_out[41]
  PIN gpio_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1161.590 0.000 1161.870 2.400 ;
    END
  END gpio_out[42]
  PIN gpio_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1409.990 0.000 1410.270 2.400 ;
    END
  END gpio_out[43]
  PIN gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 459.720 2200.000 460.320 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 557.640 2200.000 558.240 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 655.560 2200.000 656.160 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 753.480 2200.000 754.080 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 851.400 2200.000 852.000 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 949.320 2200.000 949.920 ;
    END
  END gpio_out[9]
  PIN gpio_slow_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 27.240 2200.000 27.840 ;
    END
  END gpio_slow_sel[0]
  PIN gpio_slow_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1006.440 2200.000 1007.040 ;
    END
  END gpio_slow_sel[10]
  PIN gpio_slow_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1104.360 2200.000 1104.960 ;
    END
  END gpio_slow_sel[11]
  PIN gpio_slow_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1202.280 2200.000 1202.880 ;
    END
  END gpio_slow_sel[12]
  PIN gpio_slow_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1300.200 2200.000 1300.800 ;
    END
  END gpio_slow_sel[13]
  PIN gpio_slow_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1398.120 2200.000 1398.720 ;
    END
  END gpio_slow_sel[14]
  PIN gpio_slow_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2162.090 1497.600 2162.370 1500.000 ;
    END
  END gpio_slow_sel[15]
  PIN gpio_slow_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1919.210 1497.600 1919.490 1500.000 ;
    END
  END gpio_slow_sel[16]
  PIN gpio_slow_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1676.330 1497.600 1676.610 1500.000 ;
    END
  END gpio_slow_sel[17]
  PIN gpio_slow_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1433.450 1497.600 1433.730 1500.000 ;
    END
  END gpio_slow_sel[18]
  PIN gpio_slow_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1190.570 1497.600 1190.850 1500.000 ;
    END
  END gpio_slow_sel[19]
  PIN gpio_slow_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 125.160 2200.000 125.760 ;
    END
  END gpio_slow_sel[1]
  PIN gpio_slow_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 947.690 1497.600 947.970 1500.000 ;
    END
  END gpio_slow_sel[20]
  PIN gpio_slow_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 704.810 1497.600 705.090 1500.000 ;
    END
  END gpio_slow_sel[21]
  PIN gpio_slow_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 461.930 1497.600 462.210 1500.000 ;
    END
  END gpio_slow_sel[22]
  PIN gpio_slow_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 219.050 1497.600 219.330 1500.000 ;
    END
  END gpio_slow_sel[23]
  PIN gpio_slow_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1430.760 2.400 1431.360 ;
    END
  END gpio_slow_sel[24]
  PIN gpio_slow_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 2.400 1333.440 ;
    END
  END gpio_slow_sel[25]
  PIN gpio_slow_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.920 2.400 1235.520 ;
    END
  END gpio_slow_sel[26]
  PIN gpio_slow_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 2.400 1137.600 ;
    END
  END gpio_slow_sel[27]
  PIN gpio_slow_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.080 2.400 1039.680 ;
    END
  END gpio_slow_sel[28]
  PIN gpio_slow_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 2.400 941.760 ;
    END
  END gpio_slow_sel[29]
  PIN gpio_slow_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 223.080 2200.000 223.680 ;
    END
  END gpio_slow_sel[2]
  PIN gpio_slow_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 2.400 843.840 ;
    END
  END gpio_slow_sel[30]
  PIN gpio_slow_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 2.400 745.920 ;
    END
  END gpio_slow_sel[31]
  PIN gpio_slow_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 2.400 648.000 ;
    END
  END gpio_slow_sel[32]
  PIN gpio_slow_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 2.400 550.080 ;
    END
  END gpio_slow_sel[33]
  PIN gpio_slow_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 2.400 452.160 ;
    END
  END gpio_slow_sel[34]
  PIN gpio_slow_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 2.400 354.240 ;
    END
  END gpio_slow_sel[35]
  PIN gpio_slow_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 2.400 256.320 ;
    END
  END gpio_slow_sel[36]
  PIN gpio_slow_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 2.400 158.400 ;
    END
  END gpio_slow_sel[37]
  PIN gpio_slow_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 2.400 ;
    END
  END gpio_slow_sel[38]
  PIN gpio_slow_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 2.400 ;
    END
  END gpio_slow_sel[39]
  PIN gpio_slow_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 321.000 2200.000 321.600 ;
    END
  END gpio_slow_sel[3]
  PIN gpio_slow_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 2.400 ;
    END
  END gpio_slow_sel[40]
  PIN gpio_slow_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 2.400 ;
    END
  END gpio_slow_sel[41]
  PIN gpio_slow_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 2.400 ;
    END
  END gpio_slow_sel[42]
  PIN gpio_slow_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1306.490 0.000 1306.770 2.400 ;
    END
  END gpio_slow_sel[43]
  PIN gpio_slow_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 418.920 2200.000 419.520 ;
    END
  END gpio_slow_sel[4]
  PIN gpio_slow_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 516.840 2200.000 517.440 ;
    END
  END gpio_slow_sel[5]
  PIN gpio_slow_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 614.760 2200.000 615.360 ;
    END
  END gpio_slow_sel[6]
  PIN gpio_slow_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 712.680 2200.000 713.280 ;
    END
  END gpio_slow_sel[7]
  PIN gpio_slow_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 810.600 2200.000 811.200 ;
    END
  END gpio_slow_sel[8]
  PIN gpio_slow_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 908.520 2200.000 909.120 ;
    END
  END gpio_slow_sel[9]
  PIN gpio_vtrip_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 76.200 2200.000 76.800 ;
    END
  END gpio_vtrip_sel[0]
  PIN gpio_vtrip_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1055.400 2200.000 1056.000 ;
    END
  END gpio_vtrip_sel[10]
  PIN gpio_vtrip_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1153.320 2200.000 1153.920 ;
    END
  END gpio_vtrip_sel[11]
  PIN gpio_vtrip_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1251.240 2200.000 1251.840 ;
    END
  END gpio_vtrip_sel[12]
  PIN gpio_vtrip_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1349.160 2200.000 1349.760 ;
    END
  END gpio_vtrip_sel[13]
  PIN gpio_vtrip_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 1447.080 2200.000 1447.680 ;
    END
  END gpio_vtrip_sel[14]
  PIN gpio_vtrip_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2040.650 1497.600 2040.930 1500.000 ;
    END
  END gpio_vtrip_sel[15]
  PIN gpio_vtrip_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1797.770 1497.600 1798.050 1500.000 ;
    END
  END gpio_vtrip_sel[16]
  PIN gpio_vtrip_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1554.890 1497.600 1555.170 1500.000 ;
    END
  END gpio_vtrip_sel[17]
  PIN gpio_vtrip_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1312.010 1497.600 1312.290 1500.000 ;
    END
  END gpio_vtrip_sel[18]
  PIN gpio_vtrip_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1069.130 1497.600 1069.410 1500.000 ;
    END
  END gpio_vtrip_sel[19]
  PIN gpio_vtrip_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 174.120 2200.000 174.720 ;
    END
  END gpio_vtrip_sel[1]
  PIN gpio_vtrip_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 826.250 1497.600 826.530 1500.000 ;
    END
  END gpio_vtrip_sel[20]
  PIN gpio_vtrip_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 583.370 1497.600 583.650 1500.000 ;
    END
  END gpio_vtrip_sel[21]
  PIN gpio_vtrip_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 340.490 1497.600 340.770 1500.000 ;
    END
  END gpio_vtrip_sel[22]
  PIN gpio_vtrip_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 97.610 1497.600 97.890 1500.000 ;
    END
  END gpio_vtrip_sel[23]
  PIN gpio_vtrip_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1381.800 2.400 1382.400 ;
    END
  END gpio_vtrip_sel[24]
  PIN gpio_vtrip_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1283.880 2.400 1284.480 ;
    END
  END gpio_vtrip_sel[25]
  PIN gpio_vtrip_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1185.960 2.400 1186.560 ;
    END
  END gpio_vtrip_sel[26]
  PIN gpio_vtrip_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 2.400 1088.640 ;
    END
  END gpio_vtrip_sel[27]
  PIN gpio_vtrip_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 2.400 990.720 ;
    END
  END gpio_vtrip_sel[28]
  PIN gpio_vtrip_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 2.400 892.800 ;
    END
  END gpio_vtrip_sel[29]
  PIN gpio_vtrip_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 272.040 2200.000 272.640 ;
    END
  END gpio_vtrip_sel[2]
  PIN gpio_vtrip_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 2.400 794.880 ;
    END
  END gpio_vtrip_sel[30]
  PIN gpio_vtrip_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 2.400 696.960 ;
    END
  END gpio_vtrip_sel[31]
  PIN gpio_vtrip_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 2.400 599.040 ;
    END
  END gpio_vtrip_sel[32]
  PIN gpio_vtrip_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 2.400 501.120 ;
    END
  END gpio_vtrip_sel[33]
  PIN gpio_vtrip_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 2.400 403.200 ;
    END
  END gpio_vtrip_sel[34]
  PIN gpio_vtrip_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 2.400 305.280 ;
    END
  END gpio_vtrip_sel[35]
  PIN gpio_vtrip_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 2.400 207.360 ;
    END
  END gpio_vtrip_sel[36]
  PIN gpio_vtrip_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END gpio_vtrip_sel[37]
  PIN gpio_vtrip_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 2.400 ;
    END
  END gpio_vtrip_sel[38]
  PIN gpio_vtrip_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 2.400 ;
    END
  END gpio_vtrip_sel[39]
  PIN gpio_vtrip_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 369.960 2200.000 370.560 ;
    END
  END gpio_vtrip_sel[3]
  PIN gpio_vtrip_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 2.400 ;
    END
  END gpio_vtrip_sel[40]
  PIN gpio_vtrip_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 2.400 ;
    END
  END gpio_vtrip_sel[41]
  PIN gpio_vtrip_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1182.290 0.000 1182.570 2.400 ;
    END
  END gpio_vtrip_sel[42]
  PIN gpio_vtrip_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1430.690 0.000 1430.970 2.400 ;
    END
  END gpio_vtrip_sel[43]
  PIN gpio_vtrip_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 467.880 2200.000 468.480 ;
    END
  END gpio_vtrip_sel[4]
  PIN gpio_vtrip_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 565.800 2200.000 566.400 ;
    END
  END gpio_vtrip_sel[5]
  PIN gpio_vtrip_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 663.720 2200.000 664.320 ;
    END
  END gpio_vtrip_sel[6]
  PIN gpio_vtrip_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 761.640 2200.000 762.240 ;
    END
  END gpio_vtrip_sel[7]
  PIN gpio_vtrip_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 859.560 2200.000 860.160 ;
    END
  END gpio_vtrip_sel[8]
  PIN gpio_vtrip_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2197.600 957.480 2200.000 958.080 ;
    END
  END gpio_vtrip_sel[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 2.400 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1741.190 0.000 1741.470 2.400 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1761.890 0.000 1762.170 2.400 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1782.590 0.000 1782.870 2.400 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1803.290 0.000 1803.570 2.400 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1823.990 0.000 1824.270 2.400 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1844.690 0.000 1844.970 2.400 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1865.390 0.000 1865.670 2.400 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1886.090 0.000 1886.370 2.400 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1906.790 0.000 1907.070 2.400 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1927.490 0.000 1927.770 2.400 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1554.890 0.000 1555.170 2.400 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1948.190 0.000 1948.470 2.400 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1968.890 0.000 1969.170 2.400 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1989.590 0.000 1989.870 2.400 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2010.290 0.000 2010.570 2.400 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2030.990 0.000 2031.270 2.400 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2051.690 0.000 2051.970 2.400 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2072.390 0.000 2072.670 2.400 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2093.090 0.000 2093.370 2.400 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2113.790 0.000 2114.070 2.400 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2134.490 0.000 2134.770 2.400 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1575.590 0.000 1575.870 2.400 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2155.190 0.000 2155.470 2.400 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2175.890 0.000 2176.170 2.400 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1596.290 0.000 1596.570 2.400 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1616.990 0.000 1617.270 2.400 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1637.690 0.000 1637.970 2.400 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 2.400 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1679.090 0.000 1679.370 2.400 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1699.790 0.000 1700.070 2.400 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1720.490 0.000 1720.770 2.400 ;
    END
  END mask_rev[9]
  PIN por
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END por
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 2.400 60.480 ;
    END
  END porb
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 2.400 ;
    END
  END resetb
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2194.200 1487.925 ;
      LAYER met1 ;
        RECT 0.070 9.220 2195.970 1490.520 ;
      LAYER met2 ;
        RECT 0.090 1497.320 16.370 1497.770 ;
        RECT 17.210 1497.320 36.610 1497.770 ;
        RECT 37.450 1497.320 56.850 1497.770 ;
        RECT 57.690 1497.320 77.090 1497.770 ;
        RECT 77.930 1497.320 97.330 1497.770 ;
        RECT 98.170 1497.320 117.570 1497.770 ;
        RECT 118.410 1497.320 137.810 1497.770 ;
        RECT 138.650 1497.320 158.050 1497.770 ;
        RECT 158.890 1497.320 178.290 1497.770 ;
        RECT 179.130 1497.320 198.530 1497.770 ;
        RECT 199.370 1497.320 218.770 1497.770 ;
        RECT 219.610 1497.320 239.010 1497.770 ;
        RECT 239.850 1497.320 259.250 1497.770 ;
        RECT 260.090 1497.320 279.490 1497.770 ;
        RECT 280.330 1497.320 299.730 1497.770 ;
        RECT 300.570 1497.320 319.970 1497.770 ;
        RECT 320.810 1497.320 340.210 1497.770 ;
        RECT 341.050 1497.320 360.450 1497.770 ;
        RECT 361.290 1497.320 380.690 1497.770 ;
        RECT 381.530 1497.320 400.930 1497.770 ;
        RECT 401.770 1497.320 421.170 1497.770 ;
        RECT 422.010 1497.320 441.410 1497.770 ;
        RECT 442.250 1497.320 461.650 1497.770 ;
        RECT 462.490 1497.320 481.890 1497.770 ;
        RECT 482.730 1497.320 502.130 1497.770 ;
        RECT 502.970 1497.320 522.370 1497.770 ;
        RECT 523.210 1497.320 542.610 1497.770 ;
        RECT 543.450 1497.320 562.850 1497.770 ;
        RECT 563.690 1497.320 583.090 1497.770 ;
        RECT 583.930 1497.320 603.330 1497.770 ;
        RECT 604.170 1497.320 623.570 1497.770 ;
        RECT 624.410 1497.320 643.810 1497.770 ;
        RECT 644.650 1497.320 664.050 1497.770 ;
        RECT 664.890 1497.320 684.290 1497.770 ;
        RECT 685.130 1497.320 704.530 1497.770 ;
        RECT 705.370 1497.320 724.770 1497.770 ;
        RECT 725.610 1497.320 745.010 1497.770 ;
        RECT 745.850 1497.320 765.250 1497.770 ;
        RECT 766.090 1497.320 785.490 1497.770 ;
        RECT 786.330 1497.320 805.730 1497.770 ;
        RECT 806.570 1497.320 825.970 1497.770 ;
        RECT 826.810 1497.320 846.210 1497.770 ;
        RECT 847.050 1497.320 866.450 1497.770 ;
        RECT 867.290 1497.320 886.690 1497.770 ;
        RECT 887.530 1497.320 906.930 1497.770 ;
        RECT 907.770 1497.320 927.170 1497.770 ;
        RECT 928.010 1497.320 947.410 1497.770 ;
        RECT 948.250 1497.320 967.650 1497.770 ;
        RECT 968.490 1497.320 987.890 1497.770 ;
        RECT 988.730 1497.320 1008.130 1497.770 ;
        RECT 1008.970 1497.320 1028.370 1497.770 ;
        RECT 1029.210 1497.320 1048.610 1497.770 ;
        RECT 1049.450 1497.320 1068.850 1497.770 ;
        RECT 1069.690 1497.320 1089.090 1497.770 ;
        RECT 1089.930 1497.320 1109.330 1497.770 ;
        RECT 1110.170 1497.320 1129.570 1497.770 ;
        RECT 1130.410 1497.320 1149.810 1497.770 ;
        RECT 1150.650 1497.320 1170.050 1497.770 ;
        RECT 1170.890 1497.320 1190.290 1497.770 ;
        RECT 1191.130 1497.320 1210.530 1497.770 ;
        RECT 1211.370 1497.320 1230.770 1497.770 ;
        RECT 1231.610 1497.320 1251.010 1497.770 ;
        RECT 1251.850 1497.320 1271.250 1497.770 ;
        RECT 1272.090 1497.320 1291.490 1497.770 ;
        RECT 1292.330 1497.320 1311.730 1497.770 ;
        RECT 1312.570 1497.320 1331.970 1497.770 ;
        RECT 1332.810 1497.320 1352.210 1497.770 ;
        RECT 1353.050 1497.320 1372.450 1497.770 ;
        RECT 1373.290 1497.320 1392.690 1497.770 ;
        RECT 1393.530 1497.320 1412.930 1497.770 ;
        RECT 1413.770 1497.320 1433.170 1497.770 ;
        RECT 1434.010 1497.320 1453.410 1497.770 ;
        RECT 1454.250 1497.320 1473.650 1497.770 ;
        RECT 1474.490 1497.320 1493.890 1497.770 ;
        RECT 1494.730 1497.320 1514.130 1497.770 ;
        RECT 1514.970 1497.320 1534.370 1497.770 ;
        RECT 1535.210 1497.320 1554.610 1497.770 ;
        RECT 1555.450 1497.320 1574.850 1497.770 ;
        RECT 1575.690 1497.320 1595.090 1497.770 ;
        RECT 1595.930 1497.320 1615.330 1497.770 ;
        RECT 1616.170 1497.320 1635.570 1497.770 ;
        RECT 1636.410 1497.320 1655.810 1497.770 ;
        RECT 1656.650 1497.320 1676.050 1497.770 ;
        RECT 1676.890 1497.320 1696.290 1497.770 ;
        RECT 1697.130 1497.320 1716.530 1497.770 ;
        RECT 1717.370 1497.320 1736.770 1497.770 ;
        RECT 1737.610 1497.320 1757.010 1497.770 ;
        RECT 1757.850 1497.320 1777.250 1497.770 ;
        RECT 1778.090 1497.320 1797.490 1497.770 ;
        RECT 1798.330 1497.320 1817.730 1497.770 ;
        RECT 1818.570 1497.320 1837.970 1497.770 ;
        RECT 1838.810 1497.320 1858.210 1497.770 ;
        RECT 1859.050 1497.320 1878.450 1497.770 ;
        RECT 1879.290 1497.320 1898.690 1497.770 ;
        RECT 1899.530 1497.320 1918.930 1497.770 ;
        RECT 1919.770 1497.320 1939.170 1497.770 ;
        RECT 1940.010 1497.320 1959.410 1497.770 ;
        RECT 1960.250 1497.320 1979.650 1497.770 ;
        RECT 1980.490 1497.320 1999.890 1497.770 ;
        RECT 2000.730 1497.320 2020.130 1497.770 ;
        RECT 2020.970 1497.320 2040.370 1497.770 ;
        RECT 2041.210 1497.320 2060.610 1497.770 ;
        RECT 2061.450 1497.320 2080.850 1497.770 ;
        RECT 2081.690 1497.320 2101.090 1497.770 ;
        RECT 2101.930 1497.320 2121.330 1497.770 ;
        RECT 2122.170 1497.320 2141.570 1497.770 ;
        RECT 2142.410 1497.320 2161.810 1497.770 ;
        RECT 2162.650 1497.320 2182.050 1497.770 ;
        RECT 2182.890 1497.320 2195.950 1497.770 ;
        RECT 0.090 2.680 2195.950 1497.320 ;
        RECT 0.090 1.630 22.810 2.680 ;
        RECT 23.650 1.630 43.510 2.680 ;
        RECT 44.350 1.630 64.210 2.680 ;
        RECT 65.050 1.630 84.910 2.680 ;
        RECT 85.750 1.630 105.610 2.680 ;
        RECT 106.450 1.630 126.310 2.680 ;
        RECT 127.150 1.630 147.010 2.680 ;
        RECT 147.850 1.630 167.710 2.680 ;
        RECT 168.550 1.630 188.410 2.680 ;
        RECT 189.250 1.630 209.110 2.680 ;
        RECT 209.950 1.630 229.810 2.680 ;
        RECT 230.650 1.630 250.510 2.680 ;
        RECT 251.350 1.630 271.210 2.680 ;
        RECT 272.050 1.630 291.910 2.680 ;
        RECT 292.750 1.630 312.610 2.680 ;
        RECT 313.450 1.630 333.310 2.680 ;
        RECT 334.150 1.630 354.010 2.680 ;
        RECT 354.850 1.630 374.710 2.680 ;
        RECT 375.550 1.630 395.410 2.680 ;
        RECT 396.250 1.630 416.110 2.680 ;
        RECT 416.950 1.630 436.810 2.680 ;
        RECT 437.650 1.630 457.510 2.680 ;
        RECT 458.350 1.630 478.210 2.680 ;
        RECT 479.050 1.630 498.910 2.680 ;
        RECT 499.750 1.630 519.610 2.680 ;
        RECT 520.450 1.630 540.310 2.680 ;
        RECT 541.150 1.630 561.010 2.680 ;
        RECT 561.850 1.630 581.710 2.680 ;
        RECT 582.550 1.630 602.410 2.680 ;
        RECT 603.250 1.630 623.110 2.680 ;
        RECT 623.950 1.630 643.810 2.680 ;
        RECT 644.650 1.630 664.510 2.680 ;
        RECT 665.350 1.630 685.210 2.680 ;
        RECT 686.050 1.630 705.910 2.680 ;
        RECT 706.750 1.630 726.610 2.680 ;
        RECT 727.450 1.630 747.310 2.680 ;
        RECT 748.150 1.630 768.010 2.680 ;
        RECT 768.850 1.630 788.710 2.680 ;
        RECT 789.550 1.630 809.410 2.680 ;
        RECT 810.250 1.630 830.110 2.680 ;
        RECT 830.950 1.630 850.810 2.680 ;
        RECT 851.650 1.630 871.510 2.680 ;
        RECT 872.350 1.630 892.210 2.680 ;
        RECT 893.050 1.630 912.910 2.680 ;
        RECT 913.750 1.630 933.610 2.680 ;
        RECT 934.450 1.630 954.310 2.680 ;
        RECT 955.150 1.630 975.010 2.680 ;
        RECT 975.850 1.630 995.710 2.680 ;
        RECT 996.550 1.630 1016.410 2.680 ;
        RECT 1017.250 1.630 1037.110 2.680 ;
        RECT 1037.950 1.630 1057.810 2.680 ;
        RECT 1058.650 1.630 1078.510 2.680 ;
        RECT 1079.350 1.630 1099.210 2.680 ;
        RECT 1100.050 1.630 1119.910 2.680 ;
        RECT 1120.750 1.630 1140.610 2.680 ;
        RECT 1141.450 1.630 1161.310 2.680 ;
        RECT 1162.150 1.630 1182.010 2.680 ;
        RECT 1182.850 1.630 1202.710 2.680 ;
        RECT 1203.550 1.630 1223.410 2.680 ;
        RECT 1224.250 1.630 1244.110 2.680 ;
        RECT 1244.950 1.630 1264.810 2.680 ;
        RECT 1265.650 1.630 1285.510 2.680 ;
        RECT 1286.350 1.630 1306.210 2.680 ;
        RECT 1307.050 1.630 1326.910 2.680 ;
        RECT 1327.750 1.630 1347.610 2.680 ;
        RECT 1348.450 1.630 1368.310 2.680 ;
        RECT 1369.150 1.630 1389.010 2.680 ;
        RECT 1389.850 1.630 1409.710 2.680 ;
        RECT 1410.550 1.630 1430.410 2.680 ;
        RECT 1431.250 1.630 1451.110 2.680 ;
        RECT 1451.950 1.630 1471.810 2.680 ;
        RECT 1472.650 1.630 1492.510 2.680 ;
        RECT 1493.350 1.630 1513.210 2.680 ;
        RECT 1514.050 1.630 1533.910 2.680 ;
        RECT 1534.750 1.630 1554.610 2.680 ;
        RECT 1555.450 1.630 1575.310 2.680 ;
        RECT 1576.150 1.630 1596.010 2.680 ;
        RECT 1596.850 1.630 1616.710 2.680 ;
        RECT 1617.550 1.630 1637.410 2.680 ;
        RECT 1638.250 1.630 1658.110 2.680 ;
        RECT 1658.950 1.630 1678.810 2.680 ;
        RECT 1679.650 1.630 1699.510 2.680 ;
        RECT 1700.350 1.630 1720.210 2.680 ;
        RECT 1721.050 1.630 1740.910 2.680 ;
        RECT 1741.750 1.630 1761.610 2.680 ;
        RECT 1762.450 1.630 1782.310 2.680 ;
        RECT 1783.150 1.630 1803.010 2.680 ;
        RECT 1803.850 1.630 1823.710 2.680 ;
        RECT 1824.550 1.630 1844.410 2.680 ;
        RECT 1845.250 1.630 1865.110 2.680 ;
        RECT 1865.950 1.630 1885.810 2.680 ;
        RECT 1886.650 1.630 1906.510 2.680 ;
        RECT 1907.350 1.630 1927.210 2.680 ;
        RECT 1928.050 1.630 1947.910 2.680 ;
        RECT 1948.750 1.630 1968.610 2.680 ;
        RECT 1969.450 1.630 1989.310 2.680 ;
        RECT 1990.150 1.630 2010.010 2.680 ;
        RECT 2010.850 1.630 2030.710 2.680 ;
        RECT 2031.550 1.630 2051.410 2.680 ;
        RECT 2052.250 1.630 2072.110 2.680 ;
        RECT 2072.950 1.630 2092.810 2.680 ;
        RECT 2093.650 1.630 2113.510 2.680 ;
        RECT 2114.350 1.630 2134.210 2.680 ;
        RECT 2135.050 1.630 2154.910 2.680 ;
        RECT 2155.750 1.630 2175.610 2.680 ;
        RECT 2176.450 1.630 2195.950 2.680 ;
      LAYER met3 ;
        RECT 2.400 1480.720 2197.600 1488.005 ;
        RECT 2.400 1479.320 2197.200 1480.720 ;
        RECT 2.400 1472.560 2197.600 1479.320 ;
        RECT 2.400 1471.160 2197.200 1472.560 ;
        RECT 2.400 1464.400 2197.600 1471.160 ;
        RECT 2.400 1463.000 2197.200 1464.400 ;
        RECT 2.400 1456.240 2197.600 1463.000 ;
        RECT 2.400 1454.840 2197.200 1456.240 ;
        RECT 2.400 1448.080 2197.600 1454.840 ;
        RECT 2.400 1446.680 2197.200 1448.080 ;
        RECT 2.400 1439.920 2197.600 1446.680 ;
        RECT 2.800 1438.520 2197.200 1439.920 ;
        RECT 2.400 1431.760 2197.600 1438.520 ;
        RECT 2.800 1430.360 2197.200 1431.760 ;
        RECT 2.400 1423.600 2197.600 1430.360 ;
        RECT 2.800 1422.200 2197.200 1423.600 ;
        RECT 2.400 1415.440 2197.600 1422.200 ;
        RECT 2.800 1414.040 2197.200 1415.440 ;
        RECT 2.400 1407.280 2197.600 1414.040 ;
        RECT 2.800 1405.880 2197.200 1407.280 ;
        RECT 2.400 1399.120 2197.600 1405.880 ;
        RECT 2.800 1397.720 2197.200 1399.120 ;
        RECT 2.400 1390.960 2197.600 1397.720 ;
        RECT 2.800 1389.560 2197.200 1390.960 ;
        RECT 2.400 1382.800 2197.600 1389.560 ;
        RECT 2.800 1381.400 2197.200 1382.800 ;
        RECT 2.400 1374.640 2197.600 1381.400 ;
        RECT 2.800 1373.240 2197.200 1374.640 ;
        RECT 2.400 1366.480 2197.600 1373.240 ;
        RECT 2.800 1365.080 2197.200 1366.480 ;
        RECT 2.400 1358.320 2197.600 1365.080 ;
        RECT 2.800 1356.920 2197.200 1358.320 ;
        RECT 2.400 1350.160 2197.600 1356.920 ;
        RECT 2.800 1348.760 2197.200 1350.160 ;
        RECT 2.400 1342.000 2197.600 1348.760 ;
        RECT 2.800 1340.600 2197.200 1342.000 ;
        RECT 2.400 1333.840 2197.600 1340.600 ;
        RECT 2.800 1332.440 2197.200 1333.840 ;
        RECT 2.400 1325.680 2197.600 1332.440 ;
        RECT 2.800 1324.280 2197.200 1325.680 ;
        RECT 2.400 1317.520 2197.600 1324.280 ;
        RECT 2.800 1316.120 2197.200 1317.520 ;
        RECT 2.400 1309.360 2197.600 1316.120 ;
        RECT 2.800 1307.960 2197.200 1309.360 ;
        RECT 2.400 1301.200 2197.600 1307.960 ;
        RECT 2.800 1299.800 2197.200 1301.200 ;
        RECT 2.400 1293.040 2197.600 1299.800 ;
        RECT 2.800 1291.640 2197.200 1293.040 ;
        RECT 2.400 1284.880 2197.600 1291.640 ;
        RECT 2.800 1283.480 2197.200 1284.880 ;
        RECT 2.400 1276.720 2197.600 1283.480 ;
        RECT 2.800 1275.320 2197.200 1276.720 ;
        RECT 2.400 1268.560 2197.600 1275.320 ;
        RECT 2.800 1267.160 2197.200 1268.560 ;
        RECT 2.400 1260.400 2197.600 1267.160 ;
        RECT 2.800 1259.000 2197.200 1260.400 ;
        RECT 2.400 1252.240 2197.600 1259.000 ;
        RECT 2.800 1250.840 2197.200 1252.240 ;
        RECT 2.400 1244.080 2197.600 1250.840 ;
        RECT 2.800 1242.680 2197.200 1244.080 ;
        RECT 2.400 1235.920 2197.600 1242.680 ;
        RECT 2.800 1234.520 2197.200 1235.920 ;
        RECT 2.400 1227.760 2197.600 1234.520 ;
        RECT 2.800 1226.360 2197.200 1227.760 ;
        RECT 2.400 1219.600 2197.600 1226.360 ;
        RECT 2.800 1218.200 2197.200 1219.600 ;
        RECT 2.400 1211.440 2197.600 1218.200 ;
        RECT 2.800 1210.040 2197.200 1211.440 ;
        RECT 2.400 1203.280 2197.600 1210.040 ;
        RECT 2.800 1201.880 2197.200 1203.280 ;
        RECT 2.400 1195.120 2197.600 1201.880 ;
        RECT 2.800 1193.720 2197.200 1195.120 ;
        RECT 2.400 1186.960 2197.600 1193.720 ;
        RECT 2.800 1185.560 2197.200 1186.960 ;
        RECT 2.400 1178.800 2197.600 1185.560 ;
        RECT 2.800 1177.400 2197.200 1178.800 ;
        RECT 2.400 1170.640 2197.600 1177.400 ;
        RECT 2.800 1169.240 2197.200 1170.640 ;
        RECT 2.400 1162.480 2197.600 1169.240 ;
        RECT 2.800 1161.080 2197.200 1162.480 ;
        RECT 2.400 1154.320 2197.600 1161.080 ;
        RECT 2.800 1152.920 2197.200 1154.320 ;
        RECT 2.400 1146.160 2197.600 1152.920 ;
        RECT 2.800 1144.760 2197.200 1146.160 ;
        RECT 2.400 1138.000 2197.600 1144.760 ;
        RECT 2.800 1136.600 2197.200 1138.000 ;
        RECT 2.400 1129.840 2197.600 1136.600 ;
        RECT 2.800 1128.440 2197.200 1129.840 ;
        RECT 2.400 1121.680 2197.600 1128.440 ;
        RECT 2.800 1120.280 2197.200 1121.680 ;
        RECT 2.400 1113.520 2197.600 1120.280 ;
        RECT 2.800 1112.120 2197.200 1113.520 ;
        RECT 2.400 1105.360 2197.600 1112.120 ;
        RECT 2.800 1103.960 2197.200 1105.360 ;
        RECT 2.400 1097.200 2197.600 1103.960 ;
        RECT 2.800 1095.800 2197.200 1097.200 ;
        RECT 2.400 1089.040 2197.600 1095.800 ;
        RECT 2.800 1087.640 2197.200 1089.040 ;
        RECT 2.400 1080.880 2197.600 1087.640 ;
        RECT 2.800 1079.480 2197.200 1080.880 ;
        RECT 2.400 1072.720 2197.600 1079.480 ;
        RECT 2.800 1071.320 2197.200 1072.720 ;
        RECT 2.400 1064.560 2197.600 1071.320 ;
        RECT 2.800 1063.160 2197.200 1064.560 ;
        RECT 2.400 1056.400 2197.600 1063.160 ;
        RECT 2.800 1055.000 2197.200 1056.400 ;
        RECT 2.400 1048.240 2197.600 1055.000 ;
        RECT 2.800 1046.840 2197.200 1048.240 ;
        RECT 2.400 1040.080 2197.600 1046.840 ;
        RECT 2.800 1038.680 2197.200 1040.080 ;
        RECT 2.400 1031.920 2197.600 1038.680 ;
        RECT 2.800 1030.520 2197.200 1031.920 ;
        RECT 2.400 1023.760 2197.600 1030.520 ;
        RECT 2.800 1022.360 2197.200 1023.760 ;
        RECT 2.400 1015.600 2197.600 1022.360 ;
        RECT 2.800 1014.200 2197.200 1015.600 ;
        RECT 2.400 1007.440 2197.600 1014.200 ;
        RECT 2.800 1006.040 2197.200 1007.440 ;
        RECT 2.400 999.280 2197.600 1006.040 ;
        RECT 2.800 997.880 2197.200 999.280 ;
        RECT 2.400 991.120 2197.600 997.880 ;
        RECT 2.800 989.720 2197.200 991.120 ;
        RECT 2.400 982.960 2197.600 989.720 ;
        RECT 2.800 981.560 2197.200 982.960 ;
        RECT 2.400 974.800 2197.600 981.560 ;
        RECT 2.800 973.400 2197.200 974.800 ;
        RECT 2.400 966.640 2197.600 973.400 ;
        RECT 2.800 965.240 2197.200 966.640 ;
        RECT 2.400 958.480 2197.600 965.240 ;
        RECT 2.800 957.080 2197.200 958.480 ;
        RECT 2.400 950.320 2197.600 957.080 ;
        RECT 2.800 948.920 2197.200 950.320 ;
        RECT 2.400 942.160 2197.600 948.920 ;
        RECT 2.800 940.760 2197.200 942.160 ;
        RECT 2.400 934.000 2197.600 940.760 ;
        RECT 2.800 932.600 2197.200 934.000 ;
        RECT 2.400 925.840 2197.600 932.600 ;
        RECT 2.800 924.440 2197.200 925.840 ;
        RECT 2.400 917.680 2197.600 924.440 ;
        RECT 2.800 916.280 2197.200 917.680 ;
        RECT 2.400 909.520 2197.600 916.280 ;
        RECT 2.800 908.120 2197.200 909.520 ;
        RECT 2.400 901.360 2197.600 908.120 ;
        RECT 2.800 899.960 2197.200 901.360 ;
        RECT 2.400 893.200 2197.600 899.960 ;
        RECT 2.800 891.800 2197.200 893.200 ;
        RECT 2.400 885.040 2197.600 891.800 ;
        RECT 2.800 883.640 2197.200 885.040 ;
        RECT 2.400 876.880 2197.600 883.640 ;
        RECT 2.800 875.480 2197.200 876.880 ;
        RECT 2.400 868.720 2197.600 875.480 ;
        RECT 2.800 867.320 2197.200 868.720 ;
        RECT 2.400 860.560 2197.600 867.320 ;
        RECT 2.800 859.160 2197.200 860.560 ;
        RECT 2.400 852.400 2197.600 859.160 ;
        RECT 2.800 851.000 2197.200 852.400 ;
        RECT 2.400 844.240 2197.600 851.000 ;
        RECT 2.800 842.840 2197.200 844.240 ;
        RECT 2.400 836.080 2197.600 842.840 ;
        RECT 2.800 834.680 2197.200 836.080 ;
        RECT 2.400 827.920 2197.600 834.680 ;
        RECT 2.800 826.520 2197.200 827.920 ;
        RECT 2.400 819.760 2197.600 826.520 ;
        RECT 2.800 818.360 2197.200 819.760 ;
        RECT 2.400 811.600 2197.600 818.360 ;
        RECT 2.800 810.200 2197.200 811.600 ;
        RECT 2.400 803.440 2197.600 810.200 ;
        RECT 2.800 802.040 2197.200 803.440 ;
        RECT 2.400 795.280 2197.600 802.040 ;
        RECT 2.800 793.880 2197.200 795.280 ;
        RECT 2.400 787.120 2197.600 793.880 ;
        RECT 2.800 785.720 2197.200 787.120 ;
        RECT 2.400 778.960 2197.600 785.720 ;
        RECT 2.800 777.560 2197.200 778.960 ;
        RECT 2.400 770.800 2197.600 777.560 ;
        RECT 2.800 769.400 2197.200 770.800 ;
        RECT 2.400 762.640 2197.600 769.400 ;
        RECT 2.800 761.240 2197.200 762.640 ;
        RECT 2.400 754.480 2197.600 761.240 ;
        RECT 2.800 753.080 2197.200 754.480 ;
        RECT 2.400 746.320 2197.600 753.080 ;
        RECT 2.800 744.920 2197.200 746.320 ;
        RECT 2.400 738.160 2197.600 744.920 ;
        RECT 2.800 736.760 2197.200 738.160 ;
        RECT 2.400 730.000 2197.600 736.760 ;
        RECT 2.800 728.600 2197.200 730.000 ;
        RECT 2.400 721.840 2197.600 728.600 ;
        RECT 2.800 720.440 2197.200 721.840 ;
        RECT 2.400 713.680 2197.600 720.440 ;
        RECT 2.800 712.280 2197.200 713.680 ;
        RECT 2.400 705.520 2197.600 712.280 ;
        RECT 2.800 704.120 2197.200 705.520 ;
        RECT 2.400 697.360 2197.600 704.120 ;
        RECT 2.800 695.960 2197.200 697.360 ;
        RECT 2.400 689.200 2197.600 695.960 ;
        RECT 2.800 687.800 2197.200 689.200 ;
        RECT 2.400 681.040 2197.600 687.800 ;
        RECT 2.800 679.640 2197.200 681.040 ;
        RECT 2.400 672.880 2197.600 679.640 ;
        RECT 2.800 671.480 2197.200 672.880 ;
        RECT 2.400 664.720 2197.600 671.480 ;
        RECT 2.800 663.320 2197.200 664.720 ;
        RECT 2.400 656.560 2197.600 663.320 ;
        RECT 2.800 655.160 2197.200 656.560 ;
        RECT 2.400 648.400 2197.600 655.160 ;
        RECT 2.800 647.000 2197.200 648.400 ;
        RECT 2.400 640.240 2197.600 647.000 ;
        RECT 2.800 638.840 2197.200 640.240 ;
        RECT 2.400 632.080 2197.600 638.840 ;
        RECT 2.800 630.680 2197.200 632.080 ;
        RECT 2.400 623.920 2197.600 630.680 ;
        RECT 2.800 622.520 2197.200 623.920 ;
        RECT 2.400 615.760 2197.600 622.520 ;
        RECT 2.800 614.360 2197.200 615.760 ;
        RECT 2.400 607.600 2197.600 614.360 ;
        RECT 2.800 606.200 2197.200 607.600 ;
        RECT 2.400 599.440 2197.600 606.200 ;
        RECT 2.800 598.040 2197.200 599.440 ;
        RECT 2.400 591.280 2197.600 598.040 ;
        RECT 2.800 589.880 2197.200 591.280 ;
        RECT 2.400 583.120 2197.600 589.880 ;
        RECT 2.800 581.720 2197.200 583.120 ;
        RECT 2.400 574.960 2197.600 581.720 ;
        RECT 2.800 573.560 2197.200 574.960 ;
        RECT 2.400 566.800 2197.600 573.560 ;
        RECT 2.800 565.400 2197.200 566.800 ;
        RECT 2.400 558.640 2197.600 565.400 ;
        RECT 2.800 557.240 2197.200 558.640 ;
        RECT 2.400 550.480 2197.600 557.240 ;
        RECT 2.800 549.080 2197.200 550.480 ;
        RECT 2.400 542.320 2197.600 549.080 ;
        RECT 2.800 540.920 2197.200 542.320 ;
        RECT 2.400 534.160 2197.600 540.920 ;
        RECT 2.800 532.760 2197.200 534.160 ;
        RECT 2.400 526.000 2197.600 532.760 ;
        RECT 2.800 524.600 2197.200 526.000 ;
        RECT 2.400 517.840 2197.600 524.600 ;
        RECT 2.800 516.440 2197.200 517.840 ;
        RECT 2.400 509.680 2197.600 516.440 ;
        RECT 2.800 508.280 2197.200 509.680 ;
        RECT 2.400 501.520 2197.600 508.280 ;
        RECT 2.800 500.120 2197.200 501.520 ;
        RECT 2.400 493.360 2197.600 500.120 ;
        RECT 2.800 491.960 2197.200 493.360 ;
        RECT 2.400 485.200 2197.600 491.960 ;
        RECT 2.800 483.800 2197.200 485.200 ;
        RECT 2.400 477.040 2197.600 483.800 ;
        RECT 2.800 475.640 2197.200 477.040 ;
        RECT 2.400 468.880 2197.600 475.640 ;
        RECT 2.800 467.480 2197.200 468.880 ;
        RECT 2.400 460.720 2197.600 467.480 ;
        RECT 2.800 459.320 2197.200 460.720 ;
        RECT 2.400 452.560 2197.600 459.320 ;
        RECT 2.800 451.160 2197.200 452.560 ;
        RECT 2.400 444.400 2197.600 451.160 ;
        RECT 2.800 443.000 2197.200 444.400 ;
        RECT 2.400 436.240 2197.600 443.000 ;
        RECT 2.800 434.840 2197.200 436.240 ;
        RECT 2.400 428.080 2197.600 434.840 ;
        RECT 2.800 426.680 2197.200 428.080 ;
        RECT 2.400 419.920 2197.600 426.680 ;
        RECT 2.800 418.520 2197.200 419.920 ;
        RECT 2.400 411.760 2197.600 418.520 ;
        RECT 2.800 410.360 2197.200 411.760 ;
        RECT 2.400 403.600 2197.600 410.360 ;
        RECT 2.800 402.200 2197.200 403.600 ;
        RECT 2.400 395.440 2197.600 402.200 ;
        RECT 2.800 394.040 2197.200 395.440 ;
        RECT 2.400 387.280 2197.600 394.040 ;
        RECT 2.800 385.880 2197.200 387.280 ;
        RECT 2.400 379.120 2197.600 385.880 ;
        RECT 2.800 377.720 2197.200 379.120 ;
        RECT 2.400 370.960 2197.600 377.720 ;
        RECT 2.800 369.560 2197.200 370.960 ;
        RECT 2.400 362.800 2197.600 369.560 ;
        RECT 2.800 361.400 2197.200 362.800 ;
        RECT 2.400 354.640 2197.600 361.400 ;
        RECT 2.800 353.240 2197.200 354.640 ;
        RECT 2.400 346.480 2197.600 353.240 ;
        RECT 2.800 345.080 2197.200 346.480 ;
        RECT 2.400 338.320 2197.600 345.080 ;
        RECT 2.800 336.920 2197.200 338.320 ;
        RECT 2.400 330.160 2197.600 336.920 ;
        RECT 2.800 328.760 2197.200 330.160 ;
        RECT 2.400 322.000 2197.600 328.760 ;
        RECT 2.800 320.600 2197.200 322.000 ;
        RECT 2.400 313.840 2197.600 320.600 ;
        RECT 2.800 312.440 2197.200 313.840 ;
        RECT 2.400 305.680 2197.600 312.440 ;
        RECT 2.800 304.280 2197.200 305.680 ;
        RECT 2.400 297.520 2197.600 304.280 ;
        RECT 2.800 296.120 2197.200 297.520 ;
        RECT 2.400 289.360 2197.600 296.120 ;
        RECT 2.800 287.960 2197.200 289.360 ;
        RECT 2.400 281.200 2197.600 287.960 ;
        RECT 2.800 279.800 2197.200 281.200 ;
        RECT 2.400 273.040 2197.600 279.800 ;
        RECT 2.800 271.640 2197.200 273.040 ;
        RECT 2.400 264.880 2197.600 271.640 ;
        RECT 2.800 263.480 2197.200 264.880 ;
        RECT 2.400 256.720 2197.600 263.480 ;
        RECT 2.800 255.320 2197.200 256.720 ;
        RECT 2.400 248.560 2197.600 255.320 ;
        RECT 2.800 247.160 2197.200 248.560 ;
        RECT 2.400 240.400 2197.600 247.160 ;
        RECT 2.800 239.000 2197.200 240.400 ;
        RECT 2.400 232.240 2197.600 239.000 ;
        RECT 2.800 230.840 2197.200 232.240 ;
        RECT 2.400 224.080 2197.600 230.840 ;
        RECT 2.800 222.680 2197.200 224.080 ;
        RECT 2.400 215.920 2197.600 222.680 ;
        RECT 2.800 214.520 2197.200 215.920 ;
        RECT 2.400 207.760 2197.600 214.520 ;
        RECT 2.800 206.360 2197.200 207.760 ;
        RECT 2.400 199.600 2197.600 206.360 ;
        RECT 2.800 198.200 2197.200 199.600 ;
        RECT 2.400 191.440 2197.600 198.200 ;
        RECT 2.800 190.040 2197.200 191.440 ;
        RECT 2.400 183.280 2197.600 190.040 ;
        RECT 2.800 181.880 2197.200 183.280 ;
        RECT 2.400 175.120 2197.600 181.880 ;
        RECT 2.800 173.720 2197.200 175.120 ;
        RECT 2.400 166.960 2197.600 173.720 ;
        RECT 2.800 165.560 2197.200 166.960 ;
        RECT 2.400 158.800 2197.600 165.560 ;
        RECT 2.800 157.400 2197.200 158.800 ;
        RECT 2.400 150.640 2197.600 157.400 ;
        RECT 2.800 149.240 2197.200 150.640 ;
        RECT 2.400 142.480 2197.600 149.240 ;
        RECT 2.800 141.080 2197.200 142.480 ;
        RECT 2.400 134.320 2197.600 141.080 ;
        RECT 2.800 132.920 2197.200 134.320 ;
        RECT 2.400 126.160 2197.600 132.920 ;
        RECT 2.800 124.760 2197.200 126.160 ;
        RECT 2.400 118.000 2197.600 124.760 ;
        RECT 2.800 116.600 2197.200 118.000 ;
        RECT 2.400 109.840 2197.600 116.600 ;
        RECT 2.800 108.440 2197.200 109.840 ;
        RECT 2.400 101.680 2197.600 108.440 ;
        RECT 2.800 100.280 2197.200 101.680 ;
        RECT 2.400 93.520 2197.600 100.280 ;
        RECT 2.800 92.120 2197.200 93.520 ;
        RECT 2.400 85.360 2197.600 92.120 ;
        RECT 2.800 83.960 2197.200 85.360 ;
        RECT 2.400 77.200 2197.600 83.960 ;
        RECT 2.800 75.800 2197.200 77.200 ;
        RECT 2.400 69.040 2197.600 75.800 ;
        RECT 2.800 67.640 2197.200 69.040 ;
        RECT 2.400 60.880 2197.600 67.640 ;
        RECT 2.800 59.480 2197.200 60.880 ;
        RECT 2.400 52.720 2197.600 59.480 ;
        RECT 2.400 51.320 2197.200 52.720 ;
        RECT 2.400 44.560 2197.600 51.320 ;
        RECT 2.400 43.160 2197.200 44.560 ;
        RECT 2.400 36.400 2197.600 43.160 ;
        RECT 2.400 35.000 2197.200 36.400 ;
        RECT 2.400 28.240 2197.600 35.000 ;
        RECT 2.400 26.840 2197.200 28.240 ;
        RECT 2.400 20.080 2197.600 26.840 ;
        RECT 2.400 18.680 2197.200 20.080 ;
        RECT 2.400 10.715 2197.600 18.680 ;
      LAYER met4 ;
        RECT 18.695 40.975 48.570 1473.385 ;
        RECT 52.470 40.975 53.670 1473.385 ;
        RECT 57.570 1046.220 88.570 1473.385 ;
        RECT 92.470 1046.220 93.670 1473.385 ;
        RECT 97.570 1046.220 128.570 1473.385 ;
        RECT 132.470 1046.220 133.670 1473.385 ;
        RECT 137.570 1046.220 168.570 1473.385 ;
        RECT 172.470 1046.220 173.670 1473.385 ;
        RECT 177.570 1046.220 208.570 1473.385 ;
        RECT 212.470 1046.220 213.670 1473.385 ;
        RECT 217.570 1046.220 248.570 1473.385 ;
        RECT 252.470 1046.840 253.670 1473.385 ;
        RECT 257.570 1046.840 288.570 1473.385 ;
        RECT 252.470 1046.560 288.570 1046.840 ;
        RECT 292.470 1046.560 293.670 1473.385 ;
        RECT 252.470 1046.220 293.670 1046.560 ;
        RECT 297.570 1046.560 328.570 1473.385 ;
        RECT 332.470 1046.560 333.670 1473.385 ;
        RECT 297.570 1046.220 333.670 1046.560 ;
        RECT 337.570 1046.220 368.570 1473.385 ;
        RECT 372.470 1046.220 373.670 1473.385 ;
        RECT 377.570 1046.220 408.570 1473.385 ;
        RECT 412.470 1046.220 413.670 1473.385 ;
        RECT 417.570 1046.220 448.570 1473.385 ;
        RECT 452.470 1046.840 453.670 1473.385 ;
        RECT 457.570 1046.840 488.570 1473.385 ;
        RECT 452.470 1046.220 488.570 1046.840 ;
        RECT 492.470 1046.220 493.670 1473.385 ;
        RECT 497.570 1046.560 528.570 1473.385 ;
        RECT 532.470 1046.560 533.670 1473.385 ;
        RECT 497.570 1046.220 533.670 1046.560 ;
        RECT 537.570 1046.220 568.570 1473.385 ;
        RECT 572.470 1046.220 573.670 1473.385 ;
        RECT 577.570 1046.220 608.570 1473.385 ;
        RECT 612.470 1046.840 613.670 1473.385 ;
        RECT 617.570 1046.840 648.570 1473.385 ;
        RECT 612.470 1046.220 648.570 1046.840 ;
        RECT 652.470 1046.220 653.670 1473.385 ;
        RECT 657.570 1046.560 688.570 1473.385 ;
        RECT 692.470 1046.560 693.670 1473.385 ;
        RECT 657.570 1046.220 693.670 1046.560 ;
        RECT 697.570 1046.220 728.570 1473.385 ;
        RECT 732.470 1046.220 733.670 1473.385 ;
        RECT 737.570 1046.220 768.570 1473.385 ;
        RECT 772.470 1046.220 773.670 1473.385 ;
        RECT 777.570 1046.220 808.570 1473.385 ;
        RECT 57.570 610.320 808.570 1046.220 ;
        RECT 57.570 40.975 88.570 610.320 ;
        RECT 92.470 40.975 93.670 610.320 ;
        RECT 97.570 40.975 128.570 610.320 ;
        RECT 132.470 40.975 133.670 610.320 ;
        RECT 137.570 40.975 168.570 610.320 ;
        RECT 172.470 40.975 173.670 610.320 ;
        RECT 177.570 609.920 373.670 610.320 ;
        RECT 177.570 609.700 213.670 609.920 ;
        RECT 177.570 40.975 208.570 609.700 ;
        RECT 212.470 40.975 213.670 609.700 ;
        RECT 217.570 609.700 253.670 609.920 ;
        RECT 217.570 40.975 248.570 609.700 ;
        RECT 252.470 40.975 253.670 609.700 ;
        RECT 257.570 609.700 293.670 609.920 ;
        RECT 257.570 40.975 288.570 609.700 ;
        RECT 292.470 40.975 293.670 609.700 ;
        RECT 297.570 609.700 333.670 609.920 ;
        RECT 297.570 40.975 328.570 609.700 ;
        RECT 332.470 40.975 333.670 609.700 ;
        RECT 337.570 609.700 373.670 609.920 ;
        RECT 337.570 40.975 368.570 609.700 ;
        RECT 372.470 40.975 373.670 609.700 ;
        RECT 377.570 40.975 408.570 610.320 ;
        RECT 412.470 609.920 448.570 610.320 ;
        RECT 412.470 40.975 413.670 609.920 ;
        RECT 417.570 40.975 448.570 609.920 ;
        RECT 452.470 609.920 493.670 610.320 ;
        RECT 452.470 40.975 453.670 609.920 ;
        RECT 457.570 609.700 493.670 609.920 ;
        RECT 457.570 40.975 488.570 609.700 ;
        RECT 492.470 40.975 493.670 609.700 ;
        RECT 497.570 609.700 533.670 610.320 ;
        RECT 497.570 40.975 528.570 609.700 ;
        RECT 532.470 40.975 533.670 609.700 ;
        RECT 537.570 40.975 568.570 610.320 ;
        RECT 572.470 40.975 573.670 610.320 ;
        RECT 577.570 40.975 608.570 610.320 ;
        RECT 612.470 609.920 648.570 610.320 ;
        RECT 612.470 40.975 613.670 609.920 ;
        RECT 617.570 40.975 648.570 609.920 ;
        RECT 652.470 40.975 653.670 610.320 ;
        RECT 657.570 40.975 688.570 610.320 ;
        RECT 692.470 40.975 693.670 610.320 ;
        RECT 697.570 40.975 728.570 610.320 ;
        RECT 732.470 40.975 733.670 610.320 ;
        RECT 737.570 40.975 768.570 610.320 ;
        RECT 772.470 40.975 773.670 610.320 ;
        RECT 777.570 40.975 808.570 610.320 ;
        RECT 812.470 40.975 813.670 1473.385 ;
        RECT 817.570 40.975 848.570 1473.385 ;
        RECT 852.470 40.975 853.670 1473.385 ;
        RECT 857.570 40.975 888.570 1473.385 ;
        RECT 892.470 40.975 893.670 1473.385 ;
        RECT 897.570 40.975 928.570 1473.385 ;
        RECT 932.470 40.975 933.670 1473.385 ;
        RECT 937.570 40.975 968.570 1473.385 ;
        RECT 972.470 40.975 973.670 1473.385 ;
        RECT 977.570 40.975 1008.570 1473.385 ;
        RECT 1012.470 40.975 1013.670 1473.385 ;
        RECT 1017.570 40.975 1048.570 1473.385 ;
        RECT 1052.470 40.975 1053.670 1473.385 ;
        RECT 1057.570 40.975 1088.570 1473.385 ;
        RECT 1092.470 40.975 1093.670 1473.385 ;
        RECT 1097.570 40.975 1128.570 1473.385 ;
        RECT 1132.470 40.975 1133.670 1473.385 ;
        RECT 1137.570 40.975 1168.570 1473.385 ;
        RECT 1172.470 40.975 1173.670 1473.385 ;
        RECT 1177.570 273.540 1208.570 1473.385 ;
        RECT 1212.470 273.540 1213.670 1473.385 ;
        RECT 1177.570 264.965 1213.670 273.540 ;
        RECT 1217.570 273.540 1248.570 1473.385 ;
        RECT 1252.470 273.540 1253.670 1473.385 ;
        RECT 1217.570 264.965 1253.670 273.540 ;
        RECT 1177.570 236.555 1253.670 264.965 ;
        RECT 1177.570 189.900 1213.670 236.555 ;
        RECT 1177.570 40.975 1208.570 189.900 ;
        RECT 1212.470 40.975 1213.670 189.900 ;
        RECT 1217.570 189.900 1253.670 236.555 ;
        RECT 1217.570 40.975 1248.570 189.900 ;
        RECT 1252.470 40.975 1253.670 189.900 ;
        RECT 1257.570 40.975 1288.570 1473.385 ;
        RECT 1292.470 40.975 1293.670 1473.385 ;
        RECT 1297.570 40.975 1328.570 1473.385 ;
        RECT 1332.470 40.975 1333.670 1473.385 ;
        RECT 1337.570 40.975 1368.570 1473.385 ;
        RECT 1372.470 40.975 1373.670 1473.385 ;
        RECT 1377.570 1046.220 1408.570 1473.385 ;
        RECT 1412.470 1046.220 1413.670 1473.385 ;
        RECT 1417.570 1046.220 1448.570 1473.385 ;
        RECT 1452.470 1046.220 1453.670 1473.385 ;
        RECT 1457.570 1046.220 1488.570 1473.385 ;
        RECT 1492.470 1046.220 1493.670 1473.385 ;
        RECT 1497.570 1046.220 1528.570 1473.385 ;
        RECT 1532.470 1046.220 1533.670 1473.385 ;
        RECT 1537.570 1046.220 1568.570 1473.385 ;
        RECT 1572.470 1046.220 1573.670 1473.385 ;
        RECT 1577.570 1046.220 1608.570 1473.385 ;
        RECT 1612.470 1046.840 1613.670 1473.385 ;
        RECT 1617.570 1046.840 1648.570 1473.385 ;
        RECT 1612.470 1046.220 1648.570 1046.840 ;
        RECT 1652.470 1046.840 1653.670 1473.385 ;
        RECT 1657.570 1046.840 1688.570 1473.385 ;
        RECT 1652.470 1046.560 1688.570 1046.840 ;
        RECT 1692.470 1046.560 1693.670 1473.385 ;
        RECT 1652.470 1046.220 1693.670 1046.560 ;
        RECT 1697.570 1046.560 1728.570 1473.385 ;
        RECT 1732.470 1046.560 1733.670 1473.385 ;
        RECT 1697.570 1046.220 1733.670 1046.560 ;
        RECT 1737.570 1046.220 1768.570 1473.385 ;
        RECT 1772.470 1046.220 1773.670 1473.385 ;
        RECT 1777.570 1046.220 1808.570 1473.385 ;
        RECT 1812.470 1046.840 1813.670 1473.385 ;
        RECT 1817.570 1046.840 1848.570 1473.385 ;
        RECT 1812.470 1046.220 1848.570 1046.840 ;
        RECT 1852.470 1046.840 1853.670 1473.385 ;
        RECT 1857.570 1046.840 1888.570 1473.385 ;
        RECT 1852.470 1046.560 1888.570 1046.840 ;
        RECT 1892.470 1046.560 1893.670 1473.385 ;
        RECT 1852.470 1046.220 1893.670 1046.560 ;
        RECT 1897.570 1046.560 1928.570 1473.385 ;
        RECT 1932.470 1046.560 1933.670 1473.385 ;
        RECT 1897.570 1046.220 1933.670 1046.560 ;
        RECT 1937.570 1046.220 1968.570 1473.385 ;
        RECT 1972.470 1046.220 1973.670 1473.385 ;
        RECT 1977.570 1046.220 2008.570 1473.385 ;
        RECT 2012.470 1046.220 2013.670 1473.385 ;
        RECT 2017.570 1046.220 2048.570 1473.385 ;
        RECT 2052.470 1046.840 2053.670 1473.385 ;
        RECT 2057.570 1046.840 2088.570 1473.385 ;
        RECT 2052.470 1046.220 2088.570 1046.840 ;
        RECT 2092.470 1046.220 2093.670 1473.385 ;
        RECT 1377.570 610.320 2093.670 1046.220 ;
        RECT 1377.570 40.975 1408.570 610.320 ;
        RECT 1412.470 40.975 1413.670 610.320 ;
        RECT 1417.570 40.975 1448.570 610.320 ;
        RECT 1452.470 40.975 1453.670 610.320 ;
        RECT 1457.570 609.920 1533.670 610.320 ;
        RECT 1457.570 609.700 1493.670 609.920 ;
        RECT 1457.570 40.975 1488.570 609.700 ;
        RECT 1492.470 40.975 1493.670 609.700 ;
        RECT 1497.570 609.700 1533.670 609.920 ;
        RECT 1497.570 40.975 1528.570 609.700 ;
        RECT 1532.470 40.975 1533.670 609.700 ;
        RECT 1537.570 609.700 1573.670 610.320 ;
        RECT 1537.570 40.975 1568.570 609.700 ;
        RECT 1572.470 40.975 1573.670 609.700 ;
        RECT 1577.570 609.920 1733.670 610.320 ;
        RECT 1577.570 609.700 1613.670 609.920 ;
        RECT 1577.570 40.975 1608.570 609.700 ;
        RECT 1612.470 40.975 1613.670 609.700 ;
        RECT 1617.570 609.700 1653.670 609.920 ;
        RECT 1617.570 40.975 1648.570 609.700 ;
        RECT 1652.470 40.975 1653.670 609.700 ;
        RECT 1657.570 609.700 1693.670 609.920 ;
        RECT 1657.570 40.975 1688.570 609.700 ;
        RECT 1692.470 40.975 1693.670 609.700 ;
        RECT 1697.570 609.700 1733.670 609.920 ;
        RECT 1697.570 40.975 1728.570 609.700 ;
        RECT 1732.470 40.975 1733.670 609.700 ;
        RECT 1737.570 40.975 1768.570 610.320 ;
        RECT 1772.470 40.975 1773.670 610.320 ;
        RECT 1777.570 40.975 1808.570 610.320 ;
        RECT 1812.470 609.920 1848.570 610.320 ;
        RECT 1812.470 40.975 1813.670 609.920 ;
        RECT 1817.570 40.975 1848.570 609.920 ;
        RECT 1852.470 609.920 1893.670 610.320 ;
        RECT 1852.470 40.975 1853.670 609.920 ;
        RECT 1857.570 609.700 1893.670 609.920 ;
        RECT 1857.570 40.975 1888.570 609.700 ;
        RECT 1892.470 40.975 1893.670 609.700 ;
        RECT 1897.570 609.700 1933.670 610.320 ;
        RECT 1897.570 40.975 1928.570 609.700 ;
        RECT 1932.470 40.975 1933.670 609.700 ;
        RECT 1937.570 40.975 1968.570 610.320 ;
        RECT 1972.470 40.975 1973.670 610.320 ;
        RECT 1977.570 40.975 2008.570 610.320 ;
        RECT 2012.470 609.920 2048.570 610.320 ;
        RECT 2012.470 40.975 2013.670 609.920 ;
        RECT 2017.570 40.975 2048.570 609.920 ;
        RECT 2052.470 40.975 2053.670 610.320 ;
        RECT 2057.570 40.975 2088.570 610.320 ;
        RECT 2092.470 40.975 2093.670 610.320 ;
        RECT 2097.570 40.975 2128.570 1473.385 ;
        RECT 2132.470 40.975 2133.670 1473.385 ;
        RECT 2137.570 40.975 2168.570 1473.385 ;
        RECT 2172.470 40.975 2173.670 1473.385 ;
        RECT 2177.570 40.975 2185.625 1473.385 ;
      LAYER met5 ;
        RECT 88.900 784.130 2091.500 811.700 ;
        RECT 88.900 744.130 2091.500 772.730 ;
        RECT 88.900 704.130 2091.500 732.730 ;
        RECT 88.900 664.130 2091.500 692.730 ;
        RECT 88.900 624.130 2091.500 652.730 ;
        RECT 88.900 584.130 2091.500 612.730 ;
        RECT 88.900 544.130 2091.500 572.730 ;
        RECT 88.900 504.130 2091.500 532.730 ;
        RECT 88.900 464.130 2091.500 492.730 ;
        RECT 88.900 424.130 2091.500 452.730 ;
        RECT 88.900 384.130 2091.500 412.730 ;
        RECT 88.900 344.130 2091.500 372.730 ;
        RECT 88.900 304.130 2091.500 332.730 ;
        RECT 88.900 264.130 2091.500 292.730 ;
        RECT 88.900 224.130 2091.500 252.730 ;
        RECT 88.900 208.300 2091.500 212.730 ;
  END
END picosoc
END LIBRARY

