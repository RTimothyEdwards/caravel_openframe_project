magic
tech sky130A
magscale 1 2
timestamp 1685879374
<< obsli1 >>
rect 1104 1071 18860 13617
<< obsm1 >>
rect 934 1040 18860 14340
<< metal2 >>
rect 1122 14200 1178 15000
rect 2594 14200 2650 15000
rect 4066 14200 4122 15000
rect 5538 14200 5594 15000
rect 7010 14200 7066 15000
rect 8482 14200 8538 15000
rect 9954 14200 10010 15000
rect 11426 14200 11482 15000
rect 12898 14200 12954 15000
rect 14370 14200 14426 15000
rect 15842 14200 15898 15000
rect 17314 14200 17370 15000
rect 18786 14200 18842 15000
rect 4986 0 5042 800
rect 14922 0 14978 800
<< obsm2 >>
rect 938 14144 1066 14362
rect 1234 14144 2538 14362
rect 2706 14144 4010 14362
rect 4178 14144 5482 14362
rect 5650 14144 6954 14362
rect 7122 14144 8426 14362
rect 8594 14144 9898 14362
rect 10066 14144 11370 14362
rect 11538 14144 12842 14362
rect 13010 14144 14314 14362
rect 14482 14144 15786 14362
rect 15954 14144 17258 14362
rect 17426 14144 18730 14362
rect 938 856 18840 14144
rect 938 734 4930 856
rect 5098 734 14866 856
rect 15034 734 18840 856
<< metal3 >>
rect 0 13336 800 13456
rect 19200 13336 20000 13456
rect 0 12520 800 12640
rect 0 11704 800 11824
rect 0 10888 800 11008
rect 19200 10888 20000 11008
rect 0 10072 800 10192
rect 0 9256 800 9376
rect 0 8440 800 8560
rect 19200 8440 20000 8560
rect 0 7624 800 7744
rect 0 6808 800 6928
rect 0 5992 800 6112
rect 19200 5992 20000 6112
rect 0 5176 800 5296
rect 0 4360 800 4480
rect 0 3544 800 3664
rect 19200 3544 20000 3664
rect 0 2728 800 2848
rect 0 1912 800 2032
rect 0 1096 800 1216
rect 19200 1096 20000 1216
<< obsm3 >>
rect 800 13536 19200 13633
rect 880 13256 19120 13536
rect 800 12720 19200 13256
rect 880 12440 19200 12720
rect 800 11904 19200 12440
rect 880 11624 19200 11904
rect 800 11088 19200 11624
rect 880 10808 19120 11088
rect 800 10272 19200 10808
rect 880 9992 19200 10272
rect 800 9456 19200 9992
rect 880 9176 19200 9456
rect 800 8640 19200 9176
rect 880 8360 19120 8640
rect 800 7824 19200 8360
rect 880 7544 19200 7824
rect 800 7008 19200 7544
rect 880 6728 19200 7008
rect 800 6192 19200 6728
rect 880 5912 19120 6192
rect 800 5376 19200 5912
rect 880 5096 19200 5376
rect 800 4560 19200 5096
rect 880 4280 19200 4560
rect 800 3744 19200 4280
rect 880 3464 19120 3744
rect 800 2928 19200 3464
rect 880 2648 19200 2928
rect 800 2112 19200 2648
rect 880 1832 19200 2112
rect 800 1296 19200 1832
rect 880 1055 19120 1296
<< metal4 >>
rect 4208 1040 4528 13648
rect 8208 1040 8528 13648
rect 12208 1040 12528 13648
rect 16208 1040 16528 13648
<< obsm4 >>
rect 9811 10371 10061 11933
<< labels >>
rlabel metal4 s 16208 1040 16528 13648 6 VGND
port 1 nsew ground default
rlabel metal4 s 8208 1040 8528 13648 6 VGND
port 1 nsew ground default
rlabel metal4 s 12208 1040 12528 13648 6 VPWR
port 2 nsew power default
rlabel metal4 s 4208 1040 4528 13648 6 VPWR
port 2 nsew power default
rlabel metal3 s 0 1096 800 1216 6 clockp[0]
port 3 nsew
rlabel metal3 s 0 1912 800 2032 6 clockp[1]
port 4 nsew
rlabel metal3 s 0 7624 800 7744 6 dco
port 5 nsew
rlabel metal3 s 0 2728 800 2848 6 div[0]
port 6 nsew
rlabel metal3 s 0 3544 800 3664 6 div[1]
port 7 nsew
rlabel metal3 s 0 4360 800 4480 6 div[2]
port 8 nsew
rlabel metal3 s 0 5176 800 5296 6 div[3]
port 9 nsew
rlabel metal3 s 0 5992 800 6112 6 div[4]
port 10 nsew
rlabel metal3 s 0 6808 800 6928 6 enable
port 11 nsew
rlabel metal3 s 0 8440 800 8560 6 ext_trim[0]
port 12 nsew
rlabel metal2 s 5538 14200 5594 15000 6 ext_trim[10]
port 13 nsew
rlabel metal2 s 7010 14200 7066 15000 6 ext_trim[11]
port 14 nsew
rlabel metal2 s 8482 14200 8538 15000 6 ext_trim[12]
port 15 nsew
rlabel metal2 s 9954 14200 10010 15000 6 ext_trim[13]
port 16 nsew
rlabel metal2 s 11426 14200 11482 15000 6 ext_trim[14]
port 17 nsew
rlabel metal2 s 12898 14200 12954 15000 6 ext_trim[15]
port 18 nsew
rlabel metal2 s 14370 14200 14426 15000 6 ext_trim[16]
port 19 nsew
rlabel metal2 s 15842 14200 15898 15000 6 ext_trim[17]
port 20 nsew
rlabel metal2 s 17314 14200 17370 15000 6 ext_trim[18]
port 21 nsew
rlabel metal2 s 18786 14200 18842 15000 6 ext_trim[19]
port 22 nsew
rlabel metal3 s 0 9256 800 9376 6 ext_trim[1]
port 23 nsew
rlabel metal3 s 19200 13336 20000 13456 6 ext_trim[20]
port 24 nsew
rlabel metal3 s 19200 10888 20000 11008 6 ext_trim[21]
port 25 nsew
rlabel metal3 s 19200 8440 20000 8560 6 ext_trim[22]
port 26 nsew
rlabel metal3 s 19200 5992 20000 6112 6 ext_trim[23]
port 27 nsew
rlabel metal3 s 19200 3544 20000 3664 6 ext_trim[24]
port 28 nsew
rlabel metal3 s 19200 1096 20000 1216 6 ext_trim[25]
port 29 nsew
rlabel metal3 s 0 10072 800 10192 6 ext_trim[2]
port 30 nsew
rlabel metal3 s 0 10888 800 11008 6 ext_trim[3]
port 31 nsew
rlabel metal3 s 0 11704 800 11824 6 ext_trim[4]
port 32 nsew
rlabel metal3 s 0 12520 800 12640 6 ext_trim[5]
port 33 nsew
rlabel metal3 s 0 13336 800 13456 6 ext_trim[6]
port 34 nsew
rlabel metal2 s 1122 14200 1178 15000 6 ext_trim[7]
port 35 nsew
rlabel metal2 s 2594 14200 2650 15000 6 ext_trim[8]
port 36 nsew
rlabel metal2 s 4066 14200 4122 15000 6 ext_trim[9]
port 37 nsew
rlabel metal2 s 14922 0 14978 800 6 osc
port 38 nsew
rlabel metal2 s 4986 0 5042 800 6 resetb
port 39 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 15000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1260958
string GDS_FILE /home/hosni/openframe/caravel_openframe_project/openlane/digital_locked_loop/runs/23_06_04_04_48/results/signoff/digital_locked_loop.magic.gds
string GDS_START 395388
<< end >>

