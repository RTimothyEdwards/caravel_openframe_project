VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO openframe_project_wrapper
  CLASS BLOCK ;
  FOREIGN openframe_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 3166.630 BY 4766.630 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 306.335 3168.750 306.685 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3222.335 3168.750 3222.685 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3447.335 3168.750 3447.685 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3672.335 3168.750 3672.685 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4118.335 3168.750 4118.685 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4564.335 3168.750 4564.685 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2981.980 4766.350 2982.260 4768.750 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.980 4766.350 2473.260 4768.750 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.980 4766.350 2216.260 4768.750 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.980 4766.350 1771.260 4768.750 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.980 4766.350 1262.260 4768.750 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 532.335 3168.750 532.685 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.980 4766.350 1004.260 4768.750 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.980 4766.350 747.260 4768.750 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.980 4766.350 490.260 4768.750 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.980 4766.350 233.260 4768.750 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 4622.945 0.280 4623.295 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3773.945 0.280 3774.295 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3557.945 0.280 3558.295 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3341.945 0.280 3342.295 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3125.945 0.280 3126.295 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2909.945 0.280 2910.295 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 757.335 3168.750 757.685 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2693.945 0.280 2694.295 ;
    END
  END analog_io[30]
  PIN analog_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2477.945 0.280 2478.295 ;
    END
  END analog_io[31]
  PIN analog_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1839.945 0.280 1840.295 ;
    END
  END analog_io[32]
  PIN analog_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1623.945 0.280 1624.295 ;
    END
  END analog_io[33]
  PIN analog_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1407.945 0.280 1408.295 ;
    END
  END analog_io[34]
  PIN analog_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1191.945 0.280 1192.295 ;
    END
  END analog_io[35]
  PIN analog_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 975.940 0.280 976.300 ;
    END
  END analog_io[36]
  PIN analog_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 759.940 0.280 760.300 ;
    END
  END analog_io[37]
  PIN analog_io[38]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.370 -2.120 738.650 0.280 ;
    END
  END analog_io[38]
  PIN analog_io[39]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.370 -2.120 1281.650 0.280 ;
    END
  END analog_io[39]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 983.335 3168.750 983.685 ;
    END
  END analog_io[3]
  PIN analog_io[40]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.370 -2.120 1555.650 0.280 ;
    END
  END analog_io[40]
  PIN analog_io[41]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.370 -2.120 1829.650 0.280 ;
    END
  END analog_io[41]
  PIN analog_io[42]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.370 -2.120 2103.650 0.280 ;
    END
  END analog_io[42]
  PIN analog_io[43]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2377.370 -2.120 2377.650 0.280 ;
    END
  END analog_io[43]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1208.335 3168.750 1208.685 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1433.335 3168.750 1433.685 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1659.335 3168.750 1659.685 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2545.335 3168.750 2545.685 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2771.335 3168.750 2771.685 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2996.335 3168.750 2996.685 ;
    END
  END analog_io[9]
  PIN analog_noesd_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 315.535 3168.750 315.885 ;
    END
  END analog_noesd_io[0]
  PIN analog_noesd_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3231.535 3168.750 3231.885 ;
    END
  END analog_noesd_io[10]
  PIN analog_noesd_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3456.535 3168.750 3456.885 ;
    END
  END analog_noesd_io[11]
  PIN analog_noesd_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3681.535 3168.750 3681.885 ;
    END
  END analog_noesd_io[12]
  PIN analog_noesd_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4127.535 3168.750 4127.885 ;
    END
  END analog_noesd_io[13]
  PIN analog_noesd_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4573.535 3168.750 4573.885 ;
    END
  END analog_noesd_io[14]
  PIN analog_noesd_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2972.780 4766.350 2973.060 4768.750 ;
    END
  END analog_noesd_io[15]
  PIN analog_noesd_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.780 4766.350 2464.060 4768.750 ;
    END
  END analog_noesd_io[16]
  PIN analog_noesd_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.780 4766.350 2207.060 4768.750 ;
    END
  END analog_noesd_io[17]
  PIN analog_noesd_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.780 4766.350 1762.060 4768.750 ;
    END
  END analog_noesd_io[18]
  PIN analog_noesd_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.780 4766.350 1253.060 4768.750 ;
    END
  END analog_noesd_io[19]
  PIN analog_noesd_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 541.535 3168.750 541.885 ;
    END
  END analog_noesd_io[1]
  PIN analog_noesd_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.780 4766.350 995.060 4768.750 ;
    END
  END analog_noesd_io[20]
  PIN analog_noesd_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.780 4766.350 738.060 4768.750 ;
    END
  END analog_noesd_io[21]
  PIN analog_noesd_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.780 4766.350 481.060 4768.750 ;
    END
  END analog_noesd_io[22]
  PIN analog_noesd_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.780 4766.350 224.060 4768.750 ;
    END
  END analog_noesd_io[23]
  PIN analog_noesd_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 4613.745 0.280 4614.095 ;
    END
  END analog_noesd_io[24]
  PIN analog_noesd_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3764.745 0.280 3765.095 ;
    END
  END analog_noesd_io[25]
  PIN analog_noesd_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3548.745 0.280 3549.095 ;
    END
  END analog_noesd_io[26]
  PIN analog_noesd_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3332.745 0.280 3333.095 ;
    END
  END analog_noesd_io[27]
  PIN analog_noesd_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3116.745 0.280 3117.095 ;
    END
  END analog_noesd_io[28]
  PIN analog_noesd_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2900.745 0.280 2901.095 ;
    END
  END analog_noesd_io[29]
  PIN analog_noesd_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 766.535 3168.750 766.885 ;
    END
  END analog_noesd_io[2]
  PIN analog_noesd_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2684.745 0.280 2685.095 ;
    END
  END analog_noesd_io[30]
  PIN analog_noesd_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2468.745 0.280 2469.095 ;
    END
  END analog_noesd_io[31]
  PIN analog_noesd_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1830.745 0.280 1831.095 ;
    END
  END analog_noesd_io[32]
  PIN analog_noesd_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1614.745 0.280 1615.095 ;
    END
  END analog_noesd_io[33]
  PIN analog_noesd_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1398.745 0.280 1399.095 ;
    END
  END analog_noesd_io[34]
  PIN analog_noesd_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1182.745 0.280 1183.095 ;
    END
  END analog_noesd_io[35]
  PIN analog_noesd_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 966.740 0.280 967.100 ;
    END
  END analog_noesd_io[36]
  PIN analog_noesd_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 750.740 0.280 751.100 ;
    END
  END analog_noesd_io[37]
  PIN analog_noesd_io[38]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.570 -2.120 747.850 0.280 ;
    END
  END analog_noesd_io[38]
  PIN analog_noesd_io[39]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.570 -2.120 1290.850 0.280 ;
    END
  END analog_noesd_io[39]
  PIN analog_noesd_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 992.535 3168.750 992.885 ;
    END
  END analog_noesd_io[3]
  PIN analog_noesd_io[40]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.570 -2.120 1564.850 0.280 ;
    END
  END analog_noesd_io[40]
  PIN analog_noesd_io[41]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.570 -2.120 1838.850 0.280 ;
    END
  END analog_noesd_io[41]
  PIN analog_noesd_io[42]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.570 -2.120 2112.850 0.280 ;
    END
  END analog_noesd_io[42]
  PIN analog_noesd_io[43]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.570 -2.120 2386.850 0.280 ;
    END
  END analog_noesd_io[43]
  PIN analog_noesd_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1217.535 3168.750 1217.885 ;
    END
  END analog_noesd_io[4]
  PIN analog_noesd_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1442.535 3168.750 1442.885 ;
    END
  END analog_noesd_io[5]
  PIN analog_noesd_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1668.535 3168.750 1668.885 ;
    END
  END analog_noesd_io[6]
  PIN analog_noesd_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2554.535 3168.750 2554.885 ;
    END
  END analog_noesd_io[7]
  PIN analog_noesd_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2780.535 3168.750 2780.885 ;
    END
  END analog_noesd_io[8]
  PIN analog_noesd_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3005.535 3168.750 3005.885 ;
    END
  END analog_noesd_io[9]
  PIN gpio_analog_en[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 318.295 3168.750 318.645 ;
    END
  END gpio_analog_en[0]
  PIN gpio_analog_en[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3234.295 3168.750 3234.645 ;
    END
  END gpio_analog_en[10]
  PIN gpio_analog_en[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3459.295 3168.750 3459.645 ;
    END
  END gpio_analog_en[11]
  PIN gpio_analog_en[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3684.295 3168.750 3684.645 ;
    END
  END gpio_analog_en[12]
  PIN gpio_analog_en[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4130.295 3168.750 4130.645 ;
    END
  END gpio_analog_en[13]
  PIN gpio_analog_en[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4576.295 3168.750 4576.645 ;
    END
  END gpio_analog_en[14]
  PIN gpio_analog_en[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2970.020 4766.350 2970.300 4768.750 ;
    END
  END gpio_analog_en[15]
  PIN gpio_analog_en[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2461.020 4766.350 2461.300 4768.750 ;
    END
  END gpio_analog_en[16]
  PIN gpio_analog_en[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2204.020 4766.350 2204.300 4768.750 ;
    END
  END gpio_analog_en[17]
  PIN gpio_analog_en[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1759.020 4766.350 1759.300 4768.750 ;
    END
  END gpio_analog_en[18]
  PIN gpio_analog_en[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1250.020 4766.350 1250.300 4768.750 ;
    END
  END gpio_analog_en[19]
  PIN gpio_analog_en[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 544.295 3168.750 544.645 ;
    END
  END gpio_analog_en[1]
  PIN gpio_analog_en[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 992.020 4766.350 992.300 4768.750 ;
    END
  END gpio_analog_en[20]
  PIN gpio_analog_en[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 735.020 4766.350 735.300 4768.750 ;
    END
  END gpio_analog_en[21]
  PIN gpio_analog_en[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 478.020 4766.350 478.300 4768.750 ;
    END
  END gpio_analog_en[22]
  PIN gpio_analog_en[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 221.020 4766.350 221.300 4768.750 ;
    END
  END gpio_analog_en[23]
  PIN gpio_analog_en[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4610.985 0.280 4611.335 ;
    END
  END gpio_analog_en[24]
  PIN gpio_analog_en[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3761.985 0.280 3762.335 ;
    END
  END gpio_analog_en[25]
  PIN gpio_analog_en[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3545.985 0.280 3546.335 ;
    END
  END gpio_analog_en[26]
  PIN gpio_analog_en[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3329.985 0.280 3330.335 ;
    END
  END gpio_analog_en[27]
  PIN gpio_analog_en[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3113.985 0.280 3114.335 ;
    END
  END gpio_analog_en[28]
  PIN gpio_analog_en[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2897.985 0.280 2898.335 ;
    END
  END gpio_analog_en[29]
  PIN gpio_analog_en[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 769.295 3168.750 769.645 ;
    END
  END gpio_analog_en[2]
  PIN gpio_analog_en[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2681.985 0.280 2682.335 ;
    END
  END gpio_analog_en[30]
  PIN gpio_analog_en[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2465.985 0.280 2466.335 ;
    END
  END gpio_analog_en[31]
  PIN gpio_analog_en[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1827.985 0.280 1828.335 ;
    END
  END gpio_analog_en[32]
  PIN gpio_analog_en[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1611.985 0.280 1612.335 ;
    END
  END gpio_analog_en[33]
  PIN gpio_analog_en[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1395.985 0.280 1396.335 ;
    END
  END gpio_analog_en[34]
  PIN gpio_analog_en[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1179.985 0.280 1180.335 ;
    END
  END gpio_analog_en[35]
  PIN gpio_analog_en[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 963.980 0.280 964.340 ;
    END
  END gpio_analog_en[36]
  PIN gpio_analog_en[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 747.980 0.280 748.340 ;
    END
  END gpio_analog_en[37]
  PIN gpio_analog_en[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 750.330 -2.120 750.610 0.280 ;
    END
  END gpio_analog_en[38]
  PIN gpio_analog_en[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1293.330 -2.120 1293.610 0.280 ;
    END
  END gpio_analog_en[39]
  PIN gpio_analog_en[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 995.295 3168.750 995.645 ;
    END
  END gpio_analog_en[3]
  PIN gpio_analog_en[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1567.330 -2.120 1567.610 0.280 ;
    END
  END gpio_analog_en[40]
  PIN gpio_analog_en[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1841.330 -2.120 1841.610 0.280 ;
    END
  END gpio_analog_en[41]
  PIN gpio_analog_en[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2115.330 -2.120 2115.610 0.280 ;
    END
  END gpio_analog_en[42]
  PIN gpio_analog_en[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2389.330 -2.120 2389.610 0.280 ;
    END
  END gpio_analog_en[43]
  PIN gpio_analog_en[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1220.295 3168.750 1220.645 ;
    END
  END gpio_analog_en[4]
  PIN gpio_analog_en[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1445.295 3168.750 1445.645 ;
    END
  END gpio_analog_en[5]
  PIN gpio_analog_en[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1671.295 3168.750 1671.645 ;
    END
  END gpio_analog_en[6]
  PIN gpio_analog_en[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2557.295 3168.750 2557.645 ;
    END
  END gpio_analog_en[7]
  PIN gpio_analog_en[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2783.295 3168.750 2783.645 ;
    END
  END gpio_analog_en[8]
  PIN gpio_analog_en[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3008.295 3168.750 3008.645 ;
    END
  END gpio_analog_en[9]
  PIN gpio_analog_pol[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 324.735 3168.750 325.085 ;
    END
  END gpio_analog_pol[0]
  PIN gpio_analog_pol[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3240.735 3168.750 3241.085 ;
    END
  END gpio_analog_pol[10]
  PIN gpio_analog_pol[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3465.735 3168.750 3466.085 ;
    END
  END gpio_analog_pol[11]
  PIN gpio_analog_pol[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3690.735 3168.750 3691.085 ;
    END
  END gpio_analog_pol[12]
  PIN gpio_analog_pol[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4136.735 3168.750 4137.085 ;
    END
  END gpio_analog_pol[13]
  PIN gpio_analog_pol[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4582.735 3168.750 4583.085 ;
    END
  END gpio_analog_pol[14]
  PIN gpio_analog_pol[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2963.580 4766.350 2963.860 4768.750 ;
    END
  END gpio_analog_pol[15]
  PIN gpio_analog_pol[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2454.580 4766.350 2454.860 4768.750 ;
    END
  END gpio_analog_pol[16]
  PIN gpio_analog_pol[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2197.580 4766.350 2197.860 4768.750 ;
    END
  END gpio_analog_pol[17]
  PIN gpio_analog_pol[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1752.580 4766.350 1752.860 4768.750 ;
    END
  END gpio_analog_pol[18]
  PIN gpio_analog_pol[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1243.580 4766.350 1243.860 4768.750 ;
    END
  END gpio_analog_pol[19]
  PIN gpio_analog_pol[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 550.735 3168.750 551.085 ;
    END
  END gpio_analog_pol[1]
  PIN gpio_analog_pol[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 985.580 4766.350 985.860 4768.750 ;
    END
  END gpio_analog_pol[20]
  PIN gpio_analog_pol[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 728.580 4766.350 728.860 4768.750 ;
    END
  END gpio_analog_pol[21]
  PIN gpio_analog_pol[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 471.580 4766.350 471.860 4768.750 ;
    END
  END gpio_analog_pol[22]
  PIN gpio_analog_pol[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 214.580 4766.350 214.860 4768.750 ;
    END
  END gpio_analog_pol[23]
  PIN gpio_analog_pol[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4604.545 0.280 4604.895 ;
    END
  END gpio_analog_pol[24]
  PIN gpio_analog_pol[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3755.545 0.280 3755.895 ;
    END
  END gpio_analog_pol[25]
  PIN gpio_analog_pol[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3539.545 0.280 3539.895 ;
    END
  END gpio_analog_pol[26]
  PIN gpio_analog_pol[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3323.545 0.280 3323.895 ;
    END
  END gpio_analog_pol[27]
  PIN gpio_analog_pol[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3107.545 0.280 3107.895 ;
    END
  END gpio_analog_pol[28]
  PIN gpio_analog_pol[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2891.545 0.280 2891.895 ;
    END
  END gpio_analog_pol[29]
  PIN gpio_analog_pol[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 775.735 3168.750 776.085 ;
    END
  END gpio_analog_pol[2]
  PIN gpio_analog_pol[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2675.545 0.280 2675.895 ;
    END
  END gpio_analog_pol[30]
  PIN gpio_analog_pol[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2459.545 0.280 2459.895 ;
    END
  END gpio_analog_pol[31]
  PIN gpio_analog_pol[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1821.545 0.280 1821.895 ;
    END
  END gpio_analog_pol[32]
  PIN gpio_analog_pol[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1605.545 0.280 1605.895 ;
    END
  END gpio_analog_pol[33]
  PIN gpio_analog_pol[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1389.545 0.280 1389.895 ;
    END
  END gpio_analog_pol[34]
  PIN gpio_analog_pol[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1173.545 0.280 1173.895 ;
    END
  END gpio_analog_pol[35]
  PIN gpio_analog_pol[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 957.540 0.280 957.900 ;
    END
  END gpio_analog_pol[36]
  PIN gpio_analog_pol[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 741.540 0.280 741.900 ;
    END
  END gpio_analog_pol[37]
  PIN gpio_analog_pol[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 756.770 -2.120 757.050 0.280 ;
    END
  END gpio_analog_pol[38]
  PIN gpio_analog_pol[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1299.770 -2.120 1300.050 0.280 ;
    END
  END gpio_analog_pol[39]
  PIN gpio_analog_pol[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1001.735 3168.750 1002.085 ;
    END
  END gpio_analog_pol[3]
  PIN gpio_analog_pol[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1573.770 -2.120 1574.050 0.280 ;
    END
  END gpio_analog_pol[40]
  PIN gpio_analog_pol[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1847.770 -2.120 1848.050 0.280 ;
    END
  END gpio_analog_pol[41]
  PIN gpio_analog_pol[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2121.770 -2.120 2122.050 0.280 ;
    END
  END gpio_analog_pol[42]
  PIN gpio_analog_pol[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2395.770 -2.120 2396.050 0.280 ;
    END
  END gpio_analog_pol[43]
  PIN gpio_analog_pol[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1226.735 3168.750 1227.085 ;
    END
  END gpio_analog_pol[4]
  PIN gpio_analog_pol[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1451.735 3168.750 1452.085 ;
    END
  END gpio_analog_pol[5]
  PIN gpio_analog_pol[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1677.735 3168.750 1678.085 ;
    END
  END gpio_analog_pol[6]
  PIN gpio_analog_pol[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2563.735 3168.750 2564.085 ;
    END
  END gpio_analog_pol[7]
  PIN gpio_analog_pol[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2789.735 3168.750 2790.085 ;
    END
  END gpio_analog_pol[8]
  PIN gpio_analog_pol[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3014.735 3168.750 3015.085 ;
    END
  END gpio_analog_pol[9]
  PIN gpio_analog_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 339.915 3168.750 340.265 ;
    END
  END gpio_analog_sel[0]
  PIN gpio_analog_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3255.915 3168.750 3256.265 ;
    END
  END gpio_analog_sel[10]
  PIN gpio_analog_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3480.915 3168.750 3481.265 ;
    END
  END gpio_analog_sel[11]
  PIN gpio_analog_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3705.915 3168.750 3706.265 ;
    END
  END gpio_analog_sel[12]
  PIN gpio_analog_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4151.915 3168.750 4152.265 ;
    END
  END gpio_analog_sel[13]
  PIN gpio_analog_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4597.915 3168.750 4598.265 ;
    END
  END gpio_analog_sel[14]
  PIN gpio_analog_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2948.400 4766.350 2948.680 4768.750 ;
    END
  END gpio_analog_sel[15]
  PIN gpio_analog_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2439.400 4766.350 2439.680 4768.750 ;
    END
  END gpio_analog_sel[16]
  PIN gpio_analog_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2182.400 4766.350 2182.680 4768.750 ;
    END
  END gpio_analog_sel[17]
  PIN gpio_analog_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1737.400 4766.350 1737.680 4768.750 ;
    END
  END gpio_analog_sel[18]
  PIN gpio_analog_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1228.400 4766.350 1228.680 4768.750 ;
    END
  END gpio_analog_sel[19]
  PIN gpio_analog_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 565.915 3168.750 566.265 ;
    END
  END gpio_analog_sel[1]
  PIN gpio_analog_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 970.400 4766.350 970.680 4768.750 ;
    END
  END gpio_analog_sel[20]
  PIN gpio_analog_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 713.400 4766.350 713.680 4768.750 ;
    END
  END gpio_analog_sel[21]
  PIN gpio_analog_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 456.400 4766.350 456.680 4768.750 ;
    END
  END gpio_analog_sel[22]
  PIN gpio_analog_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 199.400 4766.350 199.680 4768.750 ;
    END
  END gpio_analog_sel[23]
  PIN gpio_analog_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4589.365 0.280 4589.715 ;
    END
  END gpio_analog_sel[24]
  PIN gpio_analog_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3740.365 0.280 3740.715 ;
    END
  END gpio_analog_sel[25]
  PIN gpio_analog_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3524.365 0.280 3524.715 ;
    END
  END gpio_analog_sel[26]
  PIN gpio_analog_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3308.365 0.280 3308.715 ;
    END
  END gpio_analog_sel[27]
  PIN gpio_analog_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3092.365 0.280 3092.715 ;
    END
  END gpio_analog_sel[28]
  PIN gpio_analog_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2876.365 0.280 2876.715 ;
    END
  END gpio_analog_sel[29]
  PIN gpio_analog_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 790.915 3168.750 791.265 ;
    END
  END gpio_analog_sel[2]
  PIN gpio_analog_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2660.365 0.280 2660.715 ;
    END
  END gpio_analog_sel[30]
  PIN gpio_analog_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2444.365 0.280 2444.715 ;
    END
  END gpio_analog_sel[31]
  PIN gpio_analog_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1806.365 0.280 1806.715 ;
    END
  END gpio_analog_sel[32]
  PIN gpio_analog_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1590.365 0.280 1590.715 ;
    END
  END gpio_analog_sel[33]
  PIN gpio_analog_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1374.365 0.280 1374.715 ;
    END
  END gpio_analog_sel[34]
  PIN gpio_analog_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1158.365 0.280 1158.715 ;
    END
  END gpio_analog_sel[35]
  PIN gpio_analog_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 942.360 0.280 942.720 ;
    END
  END gpio_analog_sel[36]
  PIN gpio_analog_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 726.360 0.280 726.720 ;
    END
  END gpio_analog_sel[37]
  PIN gpio_analog_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 771.950 -2.120 772.230 0.280 ;
    END
  END gpio_analog_sel[38]
  PIN gpio_analog_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1314.950 -2.120 1315.230 0.280 ;
    END
  END gpio_analog_sel[39]
  PIN gpio_analog_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1016.915 3168.750 1017.265 ;
    END
  END gpio_analog_sel[3]
  PIN gpio_analog_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1588.950 -2.120 1589.230 0.280 ;
    END
  END gpio_analog_sel[40]
  PIN gpio_analog_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1862.950 -2.120 1863.230 0.280 ;
    END
  END gpio_analog_sel[41]
  PIN gpio_analog_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2136.950 -2.120 2137.230 0.280 ;
    END
  END gpio_analog_sel[42]
  PIN gpio_analog_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2410.950 -2.120 2411.230 0.280 ;
    END
  END gpio_analog_sel[43]
  PIN gpio_analog_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1241.915 3168.750 1242.265 ;
    END
  END gpio_analog_sel[4]
  PIN gpio_analog_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1466.915 3168.750 1467.265 ;
    END
  END gpio_analog_sel[5]
  PIN gpio_analog_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1692.915 3168.750 1693.265 ;
    END
  END gpio_analog_sel[6]
  PIN gpio_analog_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2578.915 3168.750 2579.265 ;
    END
  END gpio_analog_sel[7]
  PIN gpio_analog_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2804.915 3168.750 2805.265 ;
    END
  END gpio_analog_sel[8]
  PIN gpio_analog_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3029.915 3168.750 3030.265 ;
    END
  END gpio_analog_sel[9]
  PIN gpio_dm0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 321.515 3168.750 321.865 ;
    END
  END gpio_dm0[0]
  PIN gpio_dm0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3237.515 3168.750 3237.865 ;
    END
  END gpio_dm0[10]
  PIN gpio_dm0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3462.515 3168.750 3462.865 ;
    END
  END gpio_dm0[11]
  PIN gpio_dm0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3687.515 3168.750 3687.865 ;
    END
  END gpio_dm0[12]
  PIN gpio_dm0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4133.515 3168.750 4133.865 ;
    END
  END gpio_dm0[13]
  PIN gpio_dm0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4579.515 3168.750 4579.865 ;
    END
  END gpio_dm0[14]
  PIN gpio_dm0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2966.800 4766.350 2967.080 4768.750 ;
    END
  END gpio_dm0[15]
  PIN gpio_dm0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2457.800 4766.350 2458.080 4768.750 ;
    END
  END gpio_dm0[16]
  PIN gpio_dm0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2200.800 4766.350 2201.080 4768.750 ;
    END
  END gpio_dm0[17]
  PIN gpio_dm0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1755.800 4766.350 1756.080 4768.750 ;
    END
  END gpio_dm0[18]
  PIN gpio_dm0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1246.800 4766.350 1247.080 4768.750 ;
    END
  END gpio_dm0[19]
  PIN gpio_dm0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 547.515 3168.750 547.865 ;
    END
  END gpio_dm0[1]
  PIN gpio_dm0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 988.800 4766.350 989.080 4768.750 ;
    END
  END gpio_dm0[20]
  PIN gpio_dm0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 731.800 4766.350 732.080 4768.750 ;
    END
  END gpio_dm0[21]
  PIN gpio_dm0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 474.800 4766.350 475.080 4768.750 ;
    END
  END gpio_dm0[22]
  PIN gpio_dm0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 217.800 4766.350 218.080 4768.750 ;
    END
  END gpio_dm0[23]
  PIN gpio_dm0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4607.765 0.280 4608.115 ;
    END
  END gpio_dm0[24]
  PIN gpio_dm0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3758.765 0.280 3759.115 ;
    END
  END gpio_dm0[25]
  PIN gpio_dm0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3542.765 0.280 3543.115 ;
    END
  END gpio_dm0[26]
  PIN gpio_dm0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3326.765 0.280 3327.115 ;
    END
  END gpio_dm0[27]
  PIN gpio_dm0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3110.765 0.280 3111.115 ;
    END
  END gpio_dm0[28]
  PIN gpio_dm0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2894.765 0.280 2895.115 ;
    END
  END gpio_dm0[29]
  PIN gpio_dm0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 772.515 3168.750 772.865 ;
    END
  END gpio_dm0[2]
  PIN gpio_dm0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2678.765 0.280 2679.115 ;
    END
  END gpio_dm0[30]
  PIN gpio_dm0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2462.765 0.280 2463.115 ;
    END
  END gpio_dm0[31]
  PIN gpio_dm0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1824.765 0.280 1825.115 ;
    END
  END gpio_dm0[32]
  PIN gpio_dm0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1608.765 0.280 1609.115 ;
    END
  END gpio_dm0[33]
  PIN gpio_dm0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1392.765 0.280 1393.115 ;
    END
  END gpio_dm0[34]
  PIN gpio_dm0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1176.765 0.280 1177.115 ;
    END
  END gpio_dm0[35]
  PIN gpio_dm0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 960.760 0.280 961.120 ;
    END
  END gpio_dm0[36]
  PIN gpio_dm0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 744.760 0.280 745.120 ;
    END
  END gpio_dm0[37]
  PIN gpio_dm0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 744.350 -2.120 744.630 0.280 ;
    END
  END gpio_dm0[38]
  PIN gpio_dm0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1296.550 -2.120 1296.830 0.280 ;
    END
  END gpio_dm0[39]
  PIN gpio_dm0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 998.515 3168.750 998.865 ;
    END
  END gpio_dm0[3]
  PIN gpio_dm0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1570.550 -2.120 1570.830 0.280 ;
    END
  END gpio_dm0[40]
  PIN gpio_dm0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1844.550 -2.120 1844.830 0.280 ;
    END
  END gpio_dm0[41]
  PIN gpio_dm0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2118.550 -2.120 2118.830 0.280 ;
    END
  END gpio_dm0[42]
  PIN gpio_dm0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2392.550 -2.120 2392.830 0.280 ;
    END
  END gpio_dm0[43]
  PIN gpio_dm0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1223.515 3168.750 1223.865 ;
    END
  END gpio_dm0[4]
  PIN gpio_dm0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1448.515 3168.750 1448.865 ;
    END
  END gpio_dm0[5]
  PIN gpio_dm0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1674.515 3168.750 1674.865 ;
    END
  END gpio_dm0[6]
  PIN gpio_dm0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2560.515 3168.750 2560.865 ;
    END
  END gpio_dm0[7]
  PIN gpio_dm0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2786.515 3168.750 2786.865 ;
    END
  END gpio_dm0[8]
  PIN gpio_dm0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3011.515 3168.750 3011.865 ;
    END
  END gpio_dm0[9]
  PIN gpio_dm1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 312.315 3168.750 312.665 ;
    END
  END gpio_dm1[0]
  PIN gpio_dm1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3228.315 3168.750 3228.665 ;
    END
  END gpio_dm1[10]
  PIN gpio_dm1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3453.315 3168.750 3453.665 ;
    END
  END gpio_dm1[11]
  PIN gpio_dm1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3678.315 3168.750 3678.665 ;
    END
  END gpio_dm1[12]
  PIN gpio_dm1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4124.315 3168.750 4124.665 ;
    END
  END gpio_dm1[13]
  PIN gpio_dm1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4570.315 3168.750 4570.665 ;
    END
  END gpio_dm1[14]
  PIN gpio_dm1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2976.000 4766.350 2976.280 4768.750 ;
    END
  END gpio_dm1[15]
  PIN gpio_dm1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2467.000 4766.350 2467.280 4768.750 ;
    END
  END gpio_dm1[16]
  PIN gpio_dm1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2210.000 4766.350 2210.280 4768.750 ;
    END
  END gpio_dm1[17]
  PIN gpio_dm1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1765.000 4766.350 1765.280 4768.750 ;
    END
  END gpio_dm1[18]
  PIN gpio_dm1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1256.000 4766.350 1256.280 4768.750 ;
    END
  END gpio_dm1[19]
  PIN gpio_dm1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 538.315 3168.750 538.665 ;
    END
  END gpio_dm1[1]
  PIN gpio_dm1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 998.000 4766.350 998.280 4768.750 ;
    END
  END gpio_dm1[20]
  PIN gpio_dm1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 741.000 4766.350 741.280 4768.750 ;
    END
  END gpio_dm1[21]
  PIN gpio_dm1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 484.000 4766.350 484.280 4768.750 ;
    END
  END gpio_dm1[22]
  PIN gpio_dm1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 227.000 4766.350 227.280 4768.750 ;
    END
  END gpio_dm1[23]
  PIN gpio_dm1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4616.965 0.280 4617.315 ;
    END
  END gpio_dm1[24]
  PIN gpio_dm1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3767.965 0.280 3768.315 ;
    END
  END gpio_dm1[25]
  PIN gpio_dm1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3551.965 0.280 3552.315 ;
    END
  END gpio_dm1[26]
  PIN gpio_dm1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3335.965 0.280 3336.315 ;
    END
  END gpio_dm1[27]
  PIN gpio_dm1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3119.965 0.280 3120.315 ;
    END
  END gpio_dm1[28]
  PIN gpio_dm1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2903.965 0.280 2904.315 ;
    END
  END gpio_dm1[29]
  PIN gpio_dm1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 763.315 3168.750 763.665 ;
    END
  END gpio_dm1[2]
  PIN gpio_dm1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2687.965 0.280 2688.315 ;
    END
  END gpio_dm1[30]
  PIN gpio_dm1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2471.965 0.280 2472.315 ;
    END
  END gpio_dm1[31]
  PIN gpio_dm1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1833.965 0.280 1834.315 ;
    END
  END gpio_dm1[32]
  PIN gpio_dm1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1617.965 0.280 1618.315 ;
    END
  END gpio_dm1[33]
  PIN gpio_dm1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1401.965 0.280 1402.315 ;
    END
  END gpio_dm1[34]
  PIN gpio_dm1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1185.965 0.280 1186.315 ;
    END
  END gpio_dm1[35]
  PIN gpio_dm1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 969.960 0.280 970.320 ;
    END
  END gpio_dm1[36]
  PIN gpio_dm1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 753.960 0.280 754.320 ;
    END
  END gpio_dm1[37]
  PIN gpio_dm1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 753.550 -2.120 753.830 0.280 ;
    END
  END gpio_dm1[38]
  PIN gpio_dm1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1287.350 -2.120 1287.630 0.280 ;
    END
  END gpio_dm1[39]
  PIN gpio_dm1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 989.315 3168.750 989.665 ;
    END
  END gpio_dm1[3]
  PIN gpio_dm1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1561.350 -2.120 1561.630 0.280 ;
    END
  END gpio_dm1[40]
  PIN gpio_dm1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1835.350 -2.120 1835.630 0.280 ;
    END
  END gpio_dm1[41]
  PIN gpio_dm1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2109.350 -2.120 2109.630 0.280 ;
    END
  END gpio_dm1[42]
  PIN gpio_dm1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2383.350 -2.120 2383.630 0.280 ;
    END
  END gpio_dm1[43]
  PIN gpio_dm1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1214.315 3168.750 1214.665 ;
    END
  END gpio_dm1[4]
  PIN gpio_dm1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1439.315 3168.750 1439.665 ;
    END
  END gpio_dm1[5]
  PIN gpio_dm1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1665.315 3168.750 1665.665 ;
    END
  END gpio_dm1[6]
  PIN gpio_dm1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2551.315 3168.750 2551.665 ;
    END
  END gpio_dm1[7]
  PIN gpio_dm1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2777.315 3168.750 2777.665 ;
    END
  END gpio_dm1[8]
  PIN gpio_dm1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3002.315 3168.750 3002.665 ;
    END
  END gpio_dm1[9]
  PIN gpio_dm2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 343.135 3168.750 343.485 ;
    END
  END gpio_dm2[0]
  PIN gpio_dm2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3259.135 3168.750 3259.485 ;
    END
  END gpio_dm2[10]
  PIN gpio_dm2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3484.135 3168.750 3484.485 ;
    END
  END gpio_dm2[11]
  PIN gpio_dm2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3709.135 3168.750 3709.485 ;
    END
  END gpio_dm2[12]
  PIN gpio_dm2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4155.135 3168.750 4155.485 ;
    END
  END gpio_dm2[13]
  PIN gpio_dm2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4601.135 3168.750 4601.485 ;
    END
  END gpio_dm2[14]
  PIN gpio_dm2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2945.180 4766.350 2945.460 4768.750 ;
    END
  END gpio_dm2[15]
  PIN gpio_dm2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2436.180 4766.350 2436.460 4768.750 ;
    END
  END gpio_dm2[16]
  PIN gpio_dm2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2179.180 4766.350 2179.460 4768.750 ;
    END
  END gpio_dm2[17]
  PIN gpio_dm2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1734.180 4766.350 1734.460 4768.750 ;
    END
  END gpio_dm2[18]
  PIN gpio_dm2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1225.180 4766.350 1225.460 4768.750 ;
    END
  END gpio_dm2[19]
  PIN gpio_dm2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 569.135 3168.750 569.485 ;
    END
  END gpio_dm2[1]
  PIN gpio_dm2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 967.180 4766.350 967.460 4768.750 ;
    END
  END gpio_dm2[20]
  PIN gpio_dm2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 710.180 4766.350 710.460 4768.750 ;
    END
  END gpio_dm2[21]
  PIN gpio_dm2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 453.180 4766.350 453.460 4768.750 ;
    END
  END gpio_dm2[22]
  PIN gpio_dm2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 196.180 4766.350 196.460 4768.750 ;
    END
  END gpio_dm2[23]
  PIN gpio_dm2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4586.145 0.280 4586.495 ;
    END
  END gpio_dm2[24]
  PIN gpio_dm2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3737.145 0.280 3737.495 ;
    END
  END gpio_dm2[25]
  PIN gpio_dm2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3521.145 0.280 3521.495 ;
    END
  END gpio_dm2[26]
  PIN gpio_dm2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3305.145 0.280 3305.495 ;
    END
  END gpio_dm2[27]
  PIN gpio_dm2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3089.145 0.280 3089.495 ;
    END
  END gpio_dm2[28]
  PIN gpio_dm2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2873.145 0.280 2873.495 ;
    END
  END gpio_dm2[29]
  PIN gpio_dm2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 794.135 3168.750 794.485 ;
    END
  END gpio_dm2[2]
  PIN gpio_dm2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2657.145 0.280 2657.495 ;
    END
  END gpio_dm2[30]
  PIN gpio_dm2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2441.145 0.280 2441.495 ;
    END
  END gpio_dm2[31]
  PIN gpio_dm2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1803.145 0.280 1803.495 ;
    END
  END gpio_dm2[32]
  PIN gpio_dm2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1587.145 0.280 1587.495 ;
    END
  END gpio_dm2[33]
  PIN gpio_dm2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1371.145 0.280 1371.495 ;
    END
  END gpio_dm2[34]
  PIN gpio_dm2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1155.145 0.280 1155.495 ;
    END
  END gpio_dm2[35]
  PIN gpio_dm2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 939.140 0.280 939.500 ;
    END
  END gpio_dm2[36]
  PIN gpio_dm2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 723.140 0.280 723.500 ;
    END
  END gpio_dm2[37]
  PIN gpio_dm2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 775.170 -2.120 775.450 0.280 ;
    END
  END gpio_dm2[38]
  PIN gpio_dm2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1318.170 -2.120 1318.450 0.280 ;
    END
  END gpio_dm2[39]
  PIN gpio_dm2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1020.135 3168.750 1020.485 ;
    END
  END gpio_dm2[3]
  PIN gpio_dm2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1592.170 -2.120 1592.450 0.280 ;
    END
  END gpio_dm2[40]
  PIN gpio_dm2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1866.170 -2.120 1866.450 0.280 ;
    END
  END gpio_dm2[41]
  PIN gpio_dm2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2140.170 -2.120 2140.450 0.280 ;
    END
  END gpio_dm2[42]
  PIN gpio_dm2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2414.170 -2.120 2414.450 0.280 ;
    END
  END gpio_dm2[43]
  PIN gpio_dm2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1245.135 3168.750 1245.485 ;
    END
  END gpio_dm2[4]
  PIN gpio_dm2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1470.135 3168.750 1470.485 ;
    END
  END gpio_dm2[5]
  PIN gpio_dm2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1696.135 3168.750 1696.485 ;
    END
  END gpio_dm2[6]
  PIN gpio_dm2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2582.135 3168.750 2582.485 ;
    END
  END gpio_dm2[7]
  PIN gpio_dm2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2808.135 3168.750 2808.485 ;
    END
  END gpio_dm2[8]
  PIN gpio_dm2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3033.135 3168.750 3033.485 ;
    END
  END gpio_dm2[9]
  PIN gpio_holdover[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 346.355 3168.750 346.705 ;
    END
  END gpio_holdover[0]
  PIN gpio_holdover[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3262.355 3168.750 3262.705 ;
    END
  END gpio_holdover[10]
  PIN gpio_holdover[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3487.355 3168.750 3487.705 ;
    END
  END gpio_holdover[11]
  PIN gpio_holdover[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3712.355 3168.750 3712.705 ;
    END
  END gpio_holdover[12]
  PIN gpio_holdover[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4158.355 3168.750 4158.705 ;
    END
  END gpio_holdover[13]
  PIN gpio_holdover[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4604.355 3168.750 4604.705 ;
    END
  END gpio_holdover[14]
  PIN gpio_holdover[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2941.960 4766.350 2942.240 4768.750 ;
    END
  END gpio_holdover[15]
  PIN gpio_holdover[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2432.960 4766.350 2433.240 4768.750 ;
    END
  END gpio_holdover[16]
  PIN gpio_holdover[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2175.960 4766.350 2176.240 4768.750 ;
    END
  END gpio_holdover[17]
  PIN gpio_holdover[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1730.960 4766.350 1731.240 4768.750 ;
    END
  END gpio_holdover[18]
  PIN gpio_holdover[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1221.960 4766.350 1222.240 4768.750 ;
    END
  END gpio_holdover[19]
  PIN gpio_holdover[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 572.355 3168.750 572.705 ;
    END
  END gpio_holdover[1]
  PIN gpio_holdover[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 963.960 4766.350 964.240 4768.750 ;
    END
  END gpio_holdover[20]
  PIN gpio_holdover[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 706.960 4766.350 707.240 4768.750 ;
    END
  END gpio_holdover[21]
  PIN gpio_holdover[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 449.960 4766.350 450.240 4768.750 ;
    END
  END gpio_holdover[22]
  PIN gpio_holdover[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 192.960 4766.350 193.240 4768.750 ;
    END
  END gpio_holdover[23]
  PIN gpio_holdover[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4582.925 0.280 4583.275 ;
    END
  END gpio_holdover[24]
  PIN gpio_holdover[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3733.925 0.280 3734.275 ;
    END
  END gpio_holdover[25]
  PIN gpio_holdover[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3517.925 0.280 3518.275 ;
    END
  END gpio_holdover[26]
  PIN gpio_holdover[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3301.925 0.280 3302.275 ;
    END
  END gpio_holdover[27]
  PIN gpio_holdover[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3085.925 0.280 3086.275 ;
    END
  END gpio_holdover[28]
  PIN gpio_holdover[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2869.925 0.280 2870.275 ;
    END
  END gpio_holdover[29]
  PIN gpio_holdover[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 797.355 3168.750 797.705 ;
    END
  END gpio_holdover[2]
  PIN gpio_holdover[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2653.925 0.280 2654.275 ;
    END
  END gpio_holdover[30]
  PIN gpio_holdover[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2437.925 0.280 2438.275 ;
    END
  END gpio_holdover[31]
  PIN gpio_holdover[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1799.925 0.280 1800.275 ;
    END
  END gpio_holdover[32]
  PIN gpio_holdover[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1583.925 0.280 1584.275 ;
    END
  END gpio_holdover[33]
  PIN gpio_holdover[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1367.925 0.280 1368.275 ;
    END
  END gpio_holdover[34]
  PIN gpio_holdover[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1151.925 0.280 1152.275 ;
    END
  END gpio_holdover[35]
  PIN gpio_holdover[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 935.920 0.280 936.280 ;
    END
  END gpio_holdover[36]
  PIN gpio_holdover[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 719.920 0.280 720.280 ;
    END
  END gpio_holdover[37]
  PIN gpio_holdover[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 778.390 -2.120 778.670 0.280 ;
    END
  END gpio_holdover[38]
  PIN gpio_holdover[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1321.390 -2.120 1321.670 0.280 ;
    END
  END gpio_holdover[39]
  PIN gpio_holdover[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1023.355 3168.750 1023.705 ;
    END
  END gpio_holdover[3]
  PIN gpio_holdover[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1595.390 -2.120 1595.670 0.280 ;
    END
  END gpio_holdover[40]
  PIN gpio_holdover[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1869.390 -2.120 1869.670 0.280 ;
    END
  END gpio_holdover[41]
  PIN gpio_holdover[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2143.390 -2.120 2143.670 0.280 ;
    END
  END gpio_holdover[42]
  PIN gpio_holdover[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2417.390 -2.120 2417.670 0.280 ;
    END
  END gpio_holdover[43]
  PIN gpio_holdover[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1248.355 3168.750 1248.705 ;
    END
  END gpio_holdover[4]
  PIN gpio_holdover[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1473.355 3168.750 1473.705 ;
    END
  END gpio_holdover[5]
  PIN gpio_holdover[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1699.355 3168.750 1699.705 ;
    END
  END gpio_holdover[6]
  PIN gpio_holdover[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2585.355 3168.750 2585.705 ;
    END
  END gpio_holdover[7]
  PIN gpio_holdover[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2811.355 3168.750 2811.705 ;
    END
  END gpio_holdover[8]
  PIN gpio_holdover[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3036.355 3168.750 3036.705 ;
    END
  END gpio_holdover[9]
  PIN gpio_ib_mode_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 361.535 3168.750 361.885 ;
    END
  END gpio_ib_mode_sel[0]
  PIN gpio_ib_mode_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3277.535 3168.750 3277.885 ;
    END
  END gpio_ib_mode_sel[10]
  PIN gpio_ib_mode_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3502.535 3168.750 3502.885 ;
    END
  END gpio_ib_mode_sel[11]
  PIN gpio_ib_mode_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3727.535 3168.750 3727.885 ;
    END
  END gpio_ib_mode_sel[12]
  PIN gpio_ib_mode_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4173.535 3168.750 4173.885 ;
    END
  END gpio_ib_mode_sel[13]
  PIN gpio_ib_mode_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4619.535 3168.750 4619.885 ;
    END
  END gpio_ib_mode_sel[14]
  PIN gpio_ib_mode_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2926.780 4766.350 2927.060 4768.750 ;
    END
  END gpio_ib_mode_sel[15]
  PIN gpio_ib_mode_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2417.780 4766.350 2418.060 4768.750 ;
    END
  END gpio_ib_mode_sel[16]
  PIN gpio_ib_mode_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2160.780 4766.350 2161.060 4768.750 ;
    END
  END gpio_ib_mode_sel[17]
  PIN gpio_ib_mode_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1715.780 4766.350 1716.060 4768.750 ;
    END
  END gpio_ib_mode_sel[18]
  PIN gpio_ib_mode_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1206.780 4766.350 1207.060 4768.750 ;
    END
  END gpio_ib_mode_sel[19]
  PIN gpio_ib_mode_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 587.535 3168.750 587.885 ;
    END
  END gpio_ib_mode_sel[1]
  PIN gpio_ib_mode_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 948.780 4766.350 949.060 4768.750 ;
    END
  END gpio_ib_mode_sel[20]
  PIN gpio_ib_mode_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 691.780 4766.350 692.060 4768.750 ;
    END
  END gpio_ib_mode_sel[21]
  PIN gpio_ib_mode_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 434.780 4766.350 435.060 4768.750 ;
    END
  END gpio_ib_mode_sel[22]
  PIN gpio_ib_mode_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 177.780 4766.350 178.060 4768.750 ;
    END
  END gpio_ib_mode_sel[23]
  PIN gpio_ib_mode_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4567.745 0.280 4568.095 ;
    END
  END gpio_ib_mode_sel[24]
  PIN gpio_ib_mode_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3718.745 0.280 3719.095 ;
    END
  END gpio_ib_mode_sel[25]
  PIN gpio_ib_mode_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3502.745 0.280 3503.095 ;
    END
  END gpio_ib_mode_sel[26]
  PIN gpio_ib_mode_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3286.745 0.280 3287.095 ;
    END
  END gpio_ib_mode_sel[27]
  PIN gpio_ib_mode_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3070.745 0.280 3071.095 ;
    END
  END gpio_ib_mode_sel[28]
  PIN gpio_ib_mode_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2854.745 0.280 2855.095 ;
    END
  END gpio_ib_mode_sel[29]
  PIN gpio_ib_mode_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 812.535 3168.750 812.885 ;
    END
  END gpio_ib_mode_sel[2]
  PIN gpio_ib_mode_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2638.745 0.280 2639.095 ;
    END
  END gpio_ib_mode_sel[30]
  PIN gpio_ib_mode_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2422.745 0.280 2423.095 ;
    END
  END gpio_ib_mode_sel[31]
  PIN gpio_ib_mode_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1784.745 0.280 1785.095 ;
    END
  END gpio_ib_mode_sel[32]
  PIN gpio_ib_mode_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1568.745 0.280 1569.095 ;
    END
  END gpio_ib_mode_sel[33]
  PIN gpio_ib_mode_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1352.745 0.280 1353.095 ;
    END
  END gpio_ib_mode_sel[34]
  PIN gpio_ib_mode_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1136.745 0.280 1137.095 ;
    END
  END gpio_ib_mode_sel[35]
  PIN gpio_ib_mode_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 920.740 0.280 921.100 ;
    END
  END gpio_ib_mode_sel[36]
  PIN gpio_ib_mode_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 704.740 0.280 705.100 ;
    END
  END gpio_ib_mode_sel[37]
  PIN gpio_ib_mode_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 793.570 -2.120 793.850 0.280 ;
    END
  END gpio_ib_mode_sel[38]
  PIN gpio_ib_mode_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1336.570 -2.120 1336.850 0.280 ;
    END
  END gpio_ib_mode_sel[39]
  PIN gpio_ib_mode_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1038.535 3168.750 1038.885 ;
    END
  END gpio_ib_mode_sel[3]
  PIN gpio_ib_mode_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1610.570 -2.120 1610.850 0.280 ;
    END
  END gpio_ib_mode_sel[40]
  PIN gpio_ib_mode_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1884.570 -2.120 1884.850 0.280 ;
    END
  END gpio_ib_mode_sel[41]
  PIN gpio_ib_mode_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2158.570 -2.120 2158.850 0.280 ;
    END
  END gpio_ib_mode_sel[42]
  PIN gpio_ib_mode_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2432.570 -2.120 2432.850 0.280 ;
    END
  END gpio_ib_mode_sel[43]
  PIN gpio_ib_mode_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1263.535 3168.750 1263.885 ;
    END
  END gpio_ib_mode_sel[4]
  PIN gpio_ib_mode_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1488.535 3168.750 1488.885 ;
    END
  END gpio_ib_mode_sel[5]
  PIN gpio_ib_mode_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1714.535 3168.750 1714.885 ;
    END
  END gpio_ib_mode_sel[6]
  PIN gpio_ib_mode_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2600.535 3168.750 2600.885 ;
    END
  END gpio_ib_mode_sel[7]
  PIN gpio_ib_mode_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2826.535 3168.750 2826.885 ;
    END
  END gpio_ib_mode_sel[8]
  PIN gpio_ib_mode_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3051.535 3168.750 3051.885 ;
    END
  END gpio_ib_mode_sel[9]
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 293.915 3168.750 294.265 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3209.915 3168.750 3210.265 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3434.915 3168.750 3435.265 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3659.915 3168.750 3660.265 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4105.915 3168.750 4106.265 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4551.915 3168.750 4552.265 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2994.400 4766.350 2994.680 4768.750 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2485.400 4766.350 2485.680 4768.750 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2228.400 4766.350 2228.680 4768.750 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1783.400 4766.350 1783.680 4768.750 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1274.400 4766.350 1274.680 4768.750 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 519.915 3168.750 520.265 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1016.400 4766.350 1016.680 4768.750 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 759.400 4766.350 759.680 4768.750 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 502.400 4766.350 502.680 4768.750 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 245.400 4766.350 245.680 4768.750 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4635.365 0.280 4635.715 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3786.365 0.280 3786.715 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3570.365 0.280 3570.715 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3354.365 0.280 3354.715 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3138.365 0.280 3138.715 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2922.365 0.280 2922.715 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 744.915 3168.750 745.265 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2706.365 0.280 2706.715 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2490.365 0.280 2490.715 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1852.365 0.280 1852.715 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1636.365 0.280 1636.715 ;
    END
  END gpio_in[33]
  PIN gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1420.365 0.280 1420.715 ;
    END
  END gpio_in[34]
  PIN gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1204.365 0.280 1204.715 ;
    END
  END gpio_in[35]
  PIN gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 988.360 0.280 988.720 ;
    END
  END gpio_in[36]
  PIN gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -2.120 772.360 0.280 772.720 ;
    END
  END gpio_in[37]
  PIN gpio_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 725.950 -2.120 726.230 0.280 ;
    END
  END gpio_in[38]
  PIN gpio_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1268.950 -2.120 1269.230 0.280 ;
    END
  END gpio_in[39]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 970.915 3168.750 971.265 ;
    END
  END gpio_in[3]
  PIN gpio_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1542.950 -2.120 1543.230 0.280 ;
    END
  END gpio_in[40]
  PIN gpio_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1816.950 -2.120 1817.230 0.280 ;
    END
  END gpio_in[41]
  PIN gpio_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2090.950 -2.120 2091.230 0.280 ;
    END
  END gpio_in[42]
  PIN gpio_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2364.950 -2.120 2365.230 0.280 ;
    END
  END gpio_in[43]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1195.915 3168.750 1196.265 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1420.915 3168.750 1421.265 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1646.915 3168.750 1647.265 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2532.915 3168.750 2533.265 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2758.915 3168.750 2759.265 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2983.915 3168.750 2984.265 ;
    END
  END gpio_in[9]
  PIN gpio_in_h[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 367.515 3168.750 367.865 ;
    END
  END gpio_in_h[0]
  PIN gpio_in_h[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3283.515 3168.750 3283.865 ;
    END
  END gpio_in_h[10]
  PIN gpio_in_h[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3508.515 3168.750 3508.865 ;
    END
  END gpio_in_h[11]
  PIN gpio_in_h[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3733.515 3168.750 3733.865 ;
    END
  END gpio_in_h[12]
  PIN gpio_in_h[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4179.515 3168.750 4179.865 ;
    END
  END gpio_in_h[13]
  PIN gpio_in_h[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4625.515 3168.750 4625.865 ;
    END
  END gpio_in_h[14]
  PIN gpio_in_h[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2920.800 4766.350 2921.080 4768.750 ;
    END
  END gpio_in_h[15]
  PIN gpio_in_h[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.800 4766.350 2412.080 4768.750 ;
    END
  END gpio_in_h[16]
  PIN gpio_in_h[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.800 4766.350 2155.080 4768.750 ;
    END
  END gpio_in_h[17]
  PIN gpio_in_h[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.800 4766.350 1710.080 4768.750 ;
    END
  END gpio_in_h[18]
  PIN gpio_in_h[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.800 4766.350 1201.080 4768.750 ;
    END
  END gpio_in_h[19]
  PIN gpio_in_h[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 593.515 3168.750 593.865 ;
    END
  END gpio_in_h[1]
  PIN gpio_in_h[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.800 4766.350 943.080 4768.750 ;
    END
  END gpio_in_h[20]
  PIN gpio_in_h[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.800 4766.350 686.080 4768.750 ;
    END
  END gpio_in_h[21]
  PIN gpio_in_h[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.800 4766.350 429.080 4768.750 ;
    END
  END gpio_in_h[22]
  PIN gpio_in_h[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.800 4766.350 172.080 4768.750 ;
    END
  END gpio_in_h[23]
  PIN gpio_in_h[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 4561.765 0.280 4562.115 ;
    END
  END gpio_in_h[24]
  PIN gpio_in_h[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3712.765 0.280 3713.115 ;
    END
  END gpio_in_h[25]
  PIN gpio_in_h[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3496.765 0.280 3497.115 ;
    END
  END gpio_in_h[26]
  PIN gpio_in_h[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3280.765 0.280 3281.115 ;
    END
  END gpio_in_h[27]
  PIN gpio_in_h[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 3064.765 0.280 3065.115 ;
    END
  END gpio_in_h[28]
  PIN gpio_in_h[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2848.765 0.280 2849.115 ;
    END
  END gpio_in_h[29]
  PIN gpio_in_h[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 818.515 3168.750 818.865 ;
    END
  END gpio_in_h[2]
  PIN gpio_in_h[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2632.765 0.280 2633.115 ;
    END
  END gpio_in_h[30]
  PIN gpio_in_h[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 2416.765 0.280 2417.115 ;
    END
  END gpio_in_h[31]
  PIN gpio_in_h[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1778.765 0.280 1779.115 ;
    END
  END gpio_in_h[32]
  PIN gpio_in_h[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1562.765 0.280 1563.115 ;
    END
  END gpio_in_h[33]
  PIN gpio_in_h[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1346.765 0.280 1347.115 ;
    END
  END gpio_in_h[34]
  PIN gpio_in_h[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 1130.765 0.280 1131.115 ;
    END
  END gpio_in_h[35]
  PIN gpio_in_h[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 914.760 0.280 915.120 ;
    END
  END gpio_in_h[36]
  PIN gpio_in_h[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.120 698.760 0.280 699.120 ;
    END
  END gpio_in_h[37]
  PIN gpio_in_h[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.550 -2.120 799.830 0.280 ;
    END
  END gpio_in_h[38]
  PIN gpio_in_h[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.550 -2.120 1342.830 0.280 ;
    END
  END gpio_in_h[39]
  PIN gpio_in_h[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1044.515 3168.750 1044.865 ;
    END
  END gpio_in_h[3]
  PIN gpio_in_h[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.550 -2.120 1616.830 0.280 ;
    END
  END gpio_in_h[40]
  PIN gpio_in_h[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.550 -2.120 1890.830 0.280 ;
    END
  END gpio_in_h[41]
  PIN gpio_in_h[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.550 -2.120 2164.830 0.280 ;
    END
  END gpio_in_h[42]
  PIN gpio_in_h[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2438.550 -2.120 2438.830 0.280 ;
    END
  END gpio_in_h[43]
  PIN gpio_in_h[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1269.515 3168.750 1269.865 ;
    END
  END gpio_in_h[4]
  PIN gpio_in_h[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1494.515 3168.750 1494.865 ;
    END
  END gpio_in_h[5]
  PIN gpio_in_h[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1720.515 3168.750 1720.865 ;
    END
  END gpio_in_h[6]
  PIN gpio_in_h[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2606.515 3168.750 2606.865 ;
    END
  END gpio_in_h[7]
  PIN gpio_in_h[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2832.515 3168.750 2832.865 ;
    END
  END gpio_in_h[8]
  PIN gpio_in_h[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3057.515 3168.750 3057.865 ;
    END
  END gpio_in_h[9]
  PIN gpio_inp_dis[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 327.495 3168.750 327.845 ;
    END
  END gpio_inp_dis[0]
  PIN gpio_inp_dis[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3243.495 3168.750 3243.845 ;
    END
  END gpio_inp_dis[10]
  PIN gpio_inp_dis[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3468.495 3168.750 3468.845 ;
    END
  END gpio_inp_dis[11]
  PIN gpio_inp_dis[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3693.495 3168.750 3693.845 ;
    END
  END gpio_inp_dis[12]
  PIN gpio_inp_dis[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4139.495 3168.750 4139.845 ;
    END
  END gpio_inp_dis[13]
  PIN gpio_inp_dis[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4585.495 3168.750 4585.845 ;
    END
  END gpio_inp_dis[14]
  PIN gpio_inp_dis[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2960.820 4766.350 2961.100 4768.750 ;
    END
  END gpio_inp_dis[15]
  PIN gpio_inp_dis[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2451.820 4766.350 2452.100 4768.750 ;
    END
  END gpio_inp_dis[16]
  PIN gpio_inp_dis[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2194.820 4766.350 2195.100 4768.750 ;
    END
  END gpio_inp_dis[17]
  PIN gpio_inp_dis[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1749.820 4766.350 1750.100 4768.750 ;
    END
  END gpio_inp_dis[18]
  PIN gpio_inp_dis[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1240.820 4766.350 1241.100 4768.750 ;
    END
  END gpio_inp_dis[19]
  PIN gpio_inp_dis[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 553.495 3168.750 553.845 ;
    END
  END gpio_inp_dis[1]
  PIN gpio_inp_dis[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 982.820 4766.350 983.100 4768.750 ;
    END
  END gpio_inp_dis[20]
  PIN gpio_inp_dis[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 725.820 4766.350 726.100 4768.750 ;
    END
  END gpio_inp_dis[21]
  PIN gpio_inp_dis[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 468.820 4766.350 469.100 4768.750 ;
    END
  END gpio_inp_dis[22]
  PIN gpio_inp_dis[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 211.820 4766.350 212.100 4768.750 ;
    END
  END gpio_inp_dis[23]
  PIN gpio_inp_dis[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4601.785 0.280 4602.135 ;
    END
  END gpio_inp_dis[24]
  PIN gpio_inp_dis[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3752.785 0.280 3753.135 ;
    END
  END gpio_inp_dis[25]
  PIN gpio_inp_dis[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3536.785 0.280 3537.135 ;
    END
  END gpio_inp_dis[26]
  PIN gpio_inp_dis[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3320.785 0.280 3321.135 ;
    END
  END gpio_inp_dis[27]
  PIN gpio_inp_dis[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3104.785 0.280 3105.135 ;
    END
  END gpio_inp_dis[28]
  PIN gpio_inp_dis[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2888.785 0.280 2889.135 ;
    END
  END gpio_inp_dis[29]
  PIN gpio_inp_dis[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 778.495 3168.750 778.845 ;
    END
  END gpio_inp_dis[2]
  PIN gpio_inp_dis[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2672.785 0.280 2673.135 ;
    END
  END gpio_inp_dis[30]
  PIN gpio_inp_dis[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2456.785 0.280 2457.135 ;
    END
  END gpio_inp_dis[31]
  PIN gpio_inp_dis[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1818.785 0.280 1819.135 ;
    END
  END gpio_inp_dis[32]
  PIN gpio_inp_dis[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1602.785 0.280 1603.135 ;
    END
  END gpio_inp_dis[33]
  PIN gpio_inp_dis[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1386.785 0.280 1387.135 ;
    END
  END gpio_inp_dis[34]
  PIN gpio_inp_dis[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1170.785 0.280 1171.135 ;
    END
  END gpio_inp_dis[35]
  PIN gpio_inp_dis[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 954.780 0.280 955.140 ;
    END
  END gpio_inp_dis[36]
  PIN gpio_inp_dis[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 738.780 0.280 739.140 ;
    END
  END gpio_inp_dis[37]
  PIN gpio_inp_dis[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 759.530 -2.120 759.810 0.280 ;
    END
  END gpio_inp_dis[38]
  PIN gpio_inp_dis[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1302.530 -2.120 1302.810 0.280 ;
    END
  END gpio_inp_dis[39]
  PIN gpio_inp_dis[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1004.495 3168.750 1004.845 ;
    END
  END gpio_inp_dis[3]
  PIN gpio_inp_dis[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1576.530 -2.120 1576.810 0.280 ;
    END
  END gpio_inp_dis[40]
  PIN gpio_inp_dis[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1850.530 -2.120 1850.810 0.280 ;
    END
  END gpio_inp_dis[41]
  PIN gpio_inp_dis[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2124.530 -2.120 2124.810 0.280 ;
    END
  END gpio_inp_dis[42]
  PIN gpio_inp_dis[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2398.530 -2.120 2398.810 0.280 ;
    END
  END gpio_inp_dis[43]
  PIN gpio_inp_dis[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1229.495 3168.750 1229.845 ;
    END
  END gpio_inp_dis[4]
  PIN gpio_inp_dis[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1454.495 3168.750 1454.845 ;
    END
  END gpio_inp_dis[5]
  PIN gpio_inp_dis[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1680.495 3168.750 1680.845 ;
    END
  END gpio_inp_dis[6]
  PIN gpio_inp_dis[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2566.495 3168.750 2566.845 ;
    END
  END gpio_inp_dis[7]
  PIN gpio_inp_dis[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2792.495 3168.750 2792.845 ;
    END
  END gpio_inp_dis[8]
  PIN gpio_inp_dis[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3017.495 3168.750 3017.845 ;
    END
  END gpio_inp_dis[9]
  PIN gpio_loopback_one[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 380.025 3167.950 380.335 ;
    END
  END gpio_loopback_one[0]
  PIN gpio_loopback_one[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3290.025 3167.950 3290.335 ;
    END
  END gpio_loopback_one[10]
  PIN gpio_loopback_one[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3515.025 3167.950 3515.335 ;
    END
  END gpio_loopback_one[11]
  PIN gpio_loopback_one[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3740.025 3167.950 3740.335 ;
    END
  END gpio_loopback_one[12]
  PIN gpio_loopback_one[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4185.025 3167.950 4185.335 ;
    END
  END gpio_loopback_one[13]
  PIN gpio_loopback_one[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4635.025 3167.950 4635.335 ;
    END
  END gpio_loopback_one[14]
  PIN gpio_loopback_one[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2891.490 4766.350 2891.790 4767.950 ;
    END
  END gpio_loopback_one[15]
  PIN gpio_loopback_one[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2394.490 4766.350 2394.790 4767.950 ;
    END
  END gpio_loopback_one[16]
  PIN gpio_loopback_one[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2138.490 4766.350 2138.790 4767.950 ;
    END
  END gpio_loopback_one[17]
  PIN gpio_loopback_one[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1693.490 4766.350 1693.790 4767.950 ;
    END
  END gpio_loopback_one[18]
  PIN gpio_loopback_one[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1171.490 4766.350 1171.790 4767.950 ;
    END
  END gpio_loopback_one[19]
  PIN gpio_loopback_one[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 605.025 3167.950 605.335 ;
    END
  END gpio_loopback_one[1]
  PIN gpio_loopback_one[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 915.490 4766.350 915.790 4767.950 ;
    END
  END gpio_loopback_one[20]
  PIN gpio_loopback_one[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 659.490 4766.350 659.790 4767.950 ;
    END
  END gpio_loopback_one[21]
  PIN gpio_loopback_one[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 403.490 4766.350 403.790 4767.950 ;
    END
  END gpio_loopback_one[22]
  PIN gpio_loopback_one[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 147.490 4766.350 147.790 4767.950 ;
    END
  END gpio_loopback_one[23]
  PIN gpio_loopback_one[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 4533.220 0.280 4533.520 ;
    END
  END gpio_loopback_one[24]
  PIN gpio_loopback_one[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 3683.220 0.280 3683.520 ;
    END
  END gpio_loopback_one[25]
  PIN gpio_loopback_one[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -1.320 3468.220 0.280 3468.520 ;
    END
  END gpio_loopback_one[26]
  PIN gpio_loopback_one[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 3253.220 0.280 3253.520 ;
    END
  END gpio_loopback_one[27]
  PIN gpio_loopback_one[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 3038.220 0.280 3038.520 ;
    END
  END gpio_loopback_one[28]
  PIN gpio_loopback_one[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -1.320 2823.220 0.280 2823.520 ;
    END
  END gpio_loopback_one[29]
  PIN gpio_loopback_one[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 830.025 3167.950 830.335 ;
    END
  END gpio_loopback_one[2]
  PIN gpio_loopback_one[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 2608.220 0.280 2608.520 ;
    END
  END gpio_loopback_one[30]
  PIN gpio_loopback_one[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -1.320 2393.220 0.280 2393.520 ;
    END
  END gpio_loopback_one[31]
  PIN gpio_loopback_one[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 1748.220 0.280 1748.520 ;
    END
  END gpio_loopback_one[32]
  PIN gpio_loopback_one[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 1533.220 0.280 1533.520 ;
    END
  END gpio_loopback_one[33]
  PIN gpio_loopback_one[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 1318.220 0.280 1318.520 ;
    END
  END gpio_loopback_one[34]
  PIN gpio_loopback_one[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 1103.220 0.280 1103.520 ;
    END
  END gpio_loopback_one[35]
  PIN gpio_loopback_one[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 888.220 0.280 888.520 ;
    END
  END gpio_loopback_one[36]
  PIN gpio_loopback_one[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 673.220 0.280 673.520 ;
    END
  END gpio_loopback_one[37]
  PIN gpio_loopback_one[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 802.900 -1.300 803.160 0.280 ;
    END
  END gpio_loopback_one[38]
  PIN gpio_loopback_one[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1345.900 -1.300 1346.160 0.280 ;
    END
  END gpio_loopback_one[39]
  PIN gpio_loopback_one[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1055.025 3167.950 1055.335 ;
    END
  END gpio_loopback_one[3]
  PIN gpio_loopback_one[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1619.900 -1.300 1620.160 0.280 ;
    END
  END gpio_loopback_one[40]
  PIN gpio_loopback_one[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1893.900 -1.300 1894.160 0.280 ;
    END
  END gpio_loopback_one[41]
  PIN gpio_loopback_one[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2167.900 -1.300 2168.160 0.280 ;
    END
  END gpio_loopback_one[42]
  PIN gpio_loopback_one[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2441.900 -1.300 2442.160 0.280 ;
    END
  END gpio_loopback_one[43]
  PIN gpio_loopback_one[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1280.025 3167.950 1280.335 ;
    END
  END gpio_loopback_one[4]
  PIN gpio_loopback_one[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1505.025 3167.950 1505.335 ;
    END
  END gpio_loopback_one[5]
  PIN gpio_loopback_one[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1730.025 3167.950 1730.335 ;
    END
  END gpio_loopback_one[6]
  PIN gpio_loopback_one[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2615.025 3167.950 2615.335 ;
    END
  END gpio_loopback_one[7]
  PIN gpio_loopback_one[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2840.025 3167.950 2840.335 ;
    END
  END gpio_loopback_one[8]
  PIN gpio_loopback_one[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3065.025 3167.950 3065.335 ;
    END
  END gpio_loopback_one[9]
  PIN gpio_loopback_zero[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 390.035 3167.950 390.345 ;
    END
  END gpio_loopback_zero[0]
  PIN gpio_loopback_zero[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3300.035 3167.950 3300.345 ;
    END
  END gpio_loopback_zero[10]
  PIN gpio_loopback_zero[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3525.035 3167.950 3525.345 ;
    END
  END gpio_loopback_zero[11]
  PIN gpio_loopback_zero[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3750.035 3167.950 3750.345 ;
    END
  END gpio_loopback_zero[12]
  PIN gpio_loopback_zero[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4195.035 3167.950 4195.345 ;
    END
  END gpio_loopback_zero[13]
  PIN gpio_loopback_zero[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4645.035 3167.950 4645.345 ;
    END
  END gpio_loopback_zero[14]
  PIN gpio_loopback_zero[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2881.490 4766.350 2881.790 4767.950 ;
    END
  END gpio_loopback_zero[15]
  PIN gpio_loopback_zero[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2384.490 4766.350 2384.790 4767.950 ;
    END
  END gpio_loopback_zero[16]
  PIN gpio_loopback_zero[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2128.490 4766.350 2128.790 4767.950 ;
    END
  END gpio_loopback_zero[17]
  PIN gpio_loopback_zero[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1683.490 4766.350 1683.790 4767.950 ;
    END
  END gpio_loopback_zero[18]
  PIN gpio_loopback_zero[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1161.490 4766.350 1161.790 4767.950 ;
    END
  END gpio_loopback_zero[19]
  PIN gpio_loopback_zero[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 615.035 3167.950 615.345 ;
    END
  END gpio_loopback_zero[1]
  PIN gpio_loopback_zero[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 905.490 4766.350 905.790 4767.950 ;
    END
  END gpio_loopback_zero[20]
  PIN gpio_loopback_zero[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 649.490 4766.350 649.790 4767.950 ;
    END
  END gpio_loopback_zero[21]
  PIN gpio_loopback_zero[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 393.490 4766.350 393.790 4767.950 ;
    END
  END gpio_loopback_zero[22]
  PIN gpio_loopback_zero[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 137.490 4766.350 137.790 4767.950 ;
    END
  END gpio_loopback_zero[23]
  PIN gpio_loopback_zero[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 4523.220 0.280 4523.520 ;
    END
  END gpio_loopback_zero[24]
  PIN gpio_loopback_zero[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 3673.220 0.280 3673.520 ;
    END
  END gpio_loopback_zero[25]
  PIN gpio_loopback_zero[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 3458.220 0.280 3458.520 ;
    END
  END gpio_loopback_zero[26]
  PIN gpio_loopback_zero[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -1.320 3243.220 0.280 3243.520 ;
    END
  END gpio_loopback_zero[27]
  PIN gpio_loopback_zero[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -1.320 3028.220 0.280 3028.520 ;
    END
  END gpio_loopback_zero[28]
  PIN gpio_loopback_zero[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 2813.220 0.280 2813.520 ;
    END
  END gpio_loopback_zero[29]
  PIN gpio_loopback_zero[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 840.035 3167.950 840.345 ;
    END
  END gpio_loopback_zero[2]
  PIN gpio_loopback_zero[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -1.320 2598.220 0.280 2598.520 ;
    END
  END gpio_loopback_zero[30]
  PIN gpio_loopback_zero[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT -1.320 2383.220 0.280 2383.520 ;
    END
  END gpio_loopback_zero[31]
  PIN gpio_loopback_zero[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 1738.220 0.280 1738.520 ;
    END
  END gpio_loopback_zero[32]
  PIN gpio_loopback_zero[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 1523.220 0.280 1523.520 ;
    END
  END gpio_loopback_zero[33]
  PIN gpio_loopback_zero[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -1.320 1308.220 0.280 1308.520 ;
    END
  END gpio_loopback_zero[34]
  PIN gpio_loopback_zero[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 1093.220 0.280 1093.520 ;
    END
  END gpio_loopback_zero[35]
  PIN gpio_loopback_zero[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 878.220 0.280 878.520 ;
    END
  END gpio_loopback_zero[36]
  PIN gpio_loopback_zero[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.320 663.220 0.280 663.520 ;
    END
  END gpio_loopback_zero[37]
  PIN gpio_loopback_zero[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 818.955 -1.295 819.215 0.285 ;
    END
  END gpio_loopback_zero[38]
  PIN gpio_loopback_zero[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1366.800 -1.300 1367.060 0.280 ;
    END
  END gpio_loopback_zero[39]
  PIN gpio_loopback_zero[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1065.035 3167.950 1065.345 ;
    END
  END gpio_loopback_zero[3]
  PIN gpio_loopback_zero[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1640.825 -1.410 1641.085 0.170 ;
    END
  END gpio_loopback_zero[40]
  PIN gpio_loopback_zero[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1914.890 -1.300 1915.150 0.280 ;
    END
  END gpio_loopback_zero[41]
  PIN gpio_loopback_zero[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2188.890 -1.300 2189.150 0.280 ;
    END
  END gpio_loopback_zero[42]
  PIN gpio_loopback_zero[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2463.175 -1.300 2463.435 0.280 ;
    END
  END gpio_loopback_zero[43]
  PIN gpio_loopback_zero[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1290.035 3167.950 1290.345 ;
    END
  END gpio_loopback_zero[4]
  PIN gpio_loopback_zero[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1515.035 3167.950 1515.345 ;
    END
  END gpio_loopback_zero[5]
  PIN gpio_loopback_zero[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1740.035 3167.950 1740.345 ;
    END
  END gpio_loopback_zero[6]
  PIN gpio_loopback_zero[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2625.035 3167.950 2625.345 ;
    END
  END gpio_loopback_zero[7]
  PIN gpio_loopback_zero[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2850.035 3167.950 2850.345 ;
    END
  END gpio_loopback_zero[8]
  PIN gpio_loopback_zero[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3075.035 3167.950 3075.345 ;
    END
  END gpio_loopback_zero[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 364.755 3168.750 365.105 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3280.755 3168.750 3281.105 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3505.755 3168.750 3506.105 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3730.755 3168.750 3731.105 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4176.755 3168.750 4177.105 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4622.755 3168.750 4623.105 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2923.560 4766.350 2923.840 4768.750 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2414.560 4766.350 2414.840 4768.750 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2157.560 4766.350 2157.840 4768.750 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1712.560 4766.350 1712.840 4768.750 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1203.560 4766.350 1203.840 4768.750 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 590.755 3168.750 591.105 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 945.560 4766.350 945.840 4768.750 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 688.560 4766.350 688.840 4768.750 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 431.560 4766.350 431.840 4768.750 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 174.560 4766.350 174.840 4768.750 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4564.525 0.280 4564.875 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3715.525 0.280 3715.875 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3499.525 0.280 3499.875 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3283.525 0.280 3283.875 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3067.525 0.280 3067.875 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2851.525 0.280 2851.875 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 815.755 3168.750 816.105 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2635.525 0.280 2635.875 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2419.525 0.280 2419.875 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1781.525 0.280 1781.875 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1565.525 0.280 1565.875 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1349.525 0.280 1349.875 ;
    END
  END gpio_oeb[34]
  PIN gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1133.525 0.280 1133.875 ;
    END
  END gpio_oeb[35]
  PIN gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 917.520 0.280 917.880 ;
    END
  END gpio_oeb[36]
  PIN gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 701.520 0.280 701.880 ;
    END
  END gpio_oeb[37]
  PIN gpio_oeb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 796.790 -2.120 797.070 0.280 ;
    END
  END gpio_oeb[38]
  PIN gpio_oeb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1339.790 -2.120 1340.070 0.280 ;
    END
  END gpio_oeb[39]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1041.755 3168.750 1042.105 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1613.790 -2.120 1614.070 0.280 ;
    END
  END gpio_oeb[40]
  PIN gpio_oeb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -2.120 1888.070 0.280 ;
    END
  END gpio_oeb[41]
  PIN gpio_oeb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2161.790 -2.120 2162.070 0.280 ;
    END
  END gpio_oeb[42]
  PIN gpio_oeb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2435.790 -2.120 2436.070 0.280 ;
    END
  END gpio_oeb[43]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1266.755 3168.750 1267.105 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1491.755 3168.750 1492.105 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1717.755 3168.750 1718.105 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2603.755 3168.750 2604.105 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2829.755 3168.750 2830.105 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3054.755 3168.750 3055.105 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 349.115 3168.750 349.465 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3265.115 3168.750 3265.465 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3490.115 3168.750 3490.465 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3715.115 3168.750 3715.465 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4161.115 3168.750 4161.465 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4607.115 3168.750 4607.465 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2939.200 4766.350 2939.480 4768.750 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2430.200 4766.350 2430.480 4768.750 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2173.200 4766.350 2173.480 4768.750 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1728.200 4766.350 1728.480 4768.750 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1219.200 4766.350 1219.480 4768.750 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 575.115 3168.750 575.465 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 961.200 4766.350 961.480 4768.750 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 704.200 4766.350 704.480 4768.750 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 447.200 4766.350 447.480 4768.750 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 190.200 4766.350 190.480 4768.750 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4580.165 0.280 4580.515 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3731.165 0.280 3731.515 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3515.165 0.280 3515.515 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3299.165 0.280 3299.515 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3083.165 0.280 3083.515 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2867.165 0.280 2867.515 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 800.115 3168.750 800.465 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2651.165 0.280 2651.515 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2435.165 0.280 2435.515 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1797.165 0.280 1797.515 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1581.165 0.280 1581.515 ;
    END
  END gpio_out[33]
  PIN gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1365.165 0.280 1365.515 ;
    END
  END gpio_out[34]
  PIN gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1149.165 0.280 1149.515 ;
    END
  END gpio_out[35]
  PIN gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 933.160 0.280 933.520 ;
    END
  END gpio_out[36]
  PIN gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 717.160 0.280 717.520 ;
    END
  END gpio_out[37]
  PIN gpio_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 781.150 -2.120 781.430 0.280 ;
    END
  END gpio_out[38]
  PIN gpio_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1324.150 -2.120 1324.430 0.280 ;
    END
  END gpio_out[39]
  PIN gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1026.115 3168.750 1026.465 ;
    END
  END gpio_out[3]
  PIN gpio_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1598.150 -2.120 1598.430 0.280 ;
    END
  END gpio_out[40]
  PIN gpio_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1872.150 -2.120 1872.430 0.280 ;
    END
  END gpio_out[41]
  PIN gpio_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2146.150 -2.120 2146.430 0.280 ;
    END
  END gpio_out[42]
  PIN gpio_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2420.150 -2.120 2420.430 0.280 ;
    END
  END gpio_out[43]
  PIN gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1251.115 3168.750 1251.465 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1476.115 3168.750 1476.465 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1702.115 3168.750 1702.465 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2588.115 3168.750 2588.465 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2814.115 3168.750 2814.465 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3039.115 3168.750 3039.465 ;
    END
  END gpio_out[9]
  PIN gpio_slow_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 303.115 3168.750 303.465 ;
    END
  END gpio_slow_sel[0]
  PIN gpio_slow_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3219.115 3168.750 3219.465 ;
    END
  END gpio_slow_sel[10]
  PIN gpio_slow_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3444.115 3168.750 3444.465 ;
    END
  END gpio_slow_sel[11]
  PIN gpio_slow_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3669.115 3168.750 3669.465 ;
    END
  END gpio_slow_sel[12]
  PIN gpio_slow_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4115.115 3168.750 4115.465 ;
    END
  END gpio_slow_sel[13]
  PIN gpio_slow_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4561.115 3168.750 4561.465 ;
    END
  END gpio_slow_sel[14]
  PIN gpio_slow_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2985.200 4766.350 2985.480 4768.750 ;
    END
  END gpio_slow_sel[15]
  PIN gpio_slow_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2476.200 4766.350 2476.480 4768.750 ;
    END
  END gpio_slow_sel[16]
  PIN gpio_slow_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2219.200 4766.350 2219.480 4768.750 ;
    END
  END gpio_slow_sel[17]
  PIN gpio_slow_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1774.200 4766.350 1774.480 4768.750 ;
    END
  END gpio_slow_sel[18]
  PIN gpio_slow_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1265.200 4766.350 1265.480 4768.750 ;
    END
  END gpio_slow_sel[19]
  PIN gpio_slow_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 529.115 3168.750 529.465 ;
    END
  END gpio_slow_sel[1]
  PIN gpio_slow_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1007.200 4766.350 1007.480 4768.750 ;
    END
  END gpio_slow_sel[20]
  PIN gpio_slow_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 750.200 4766.350 750.480 4768.750 ;
    END
  END gpio_slow_sel[21]
  PIN gpio_slow_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 493.200 4766.350 493.480 4768.750 ;
    END
  END gpio_slow_sel[22]
  PIN gpio_slow_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 236.200 4766.350 236.480 4768.750 ;
    END
  END gpio_slow_sel[23]
  PIN gpio_slow_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4626.165 0.280 4626.515 ;
    END
  END gpio_slow_sel[24]
  PIN gpio_slow_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3777.165 0.280 3777.515 ;
    END
  END gpio_slow_sel[25]
  PIN gpio_slow_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3561.165 0.280 3561.515 ;
    END
  END gpio_slow_sel[26]
  PIN gpio_slow_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3345.165 0.280 3345.515 ;
    END
  END gpio_slow_sel[27]
  PIN gpio_slow_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3129.165 0.280 3129.515 ;
    END
  END gpio_slow_sel[28]
  PIN gpio_slow_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2913.165 0.280 2913.515 ;
    END
  END gpio_slow_sel[29]
  PIN gpio_slow_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 754.115 3168.750 754.465 ;
    END
  END gpio_slow_sel[2]
  PIN gpio_slow_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2697.165 0.280 2697.515 ;
    END
  END gpio_slow_sel[30]
  PIN gpio_slow_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2481.165 0.280 2481.515 ;
    END
  END gpio_slow_sel[31]
  PIN gpio_slow_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1843.165 0.280 1843.515 ;
    END
  END gpio_slow_sel[32]
  PIN gpio_slow_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1627.165 0.280 1627.515 ;
    END
  END gpio_slow_sel[33]
  PIN gpio_slow_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1411.165 0.280 1411.515 ;
    END
  END gpio_slow_sel[34]
  PIN gpio_slow_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1195.165 0.280 1195.515 ;
    END
  END gpio_slow_sel[35]
  PIN gpio_slow_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 979.160 0.280 979.520 ;
    END
  END gpio_slow_sel[36]
  PIN gpio_slow_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 763.160 0.280 763.520 ;
    END
  END gpio_slow_sel[37]
  PIN gpio_slow_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 735.150 -2.120 735.430 0.280 ;
    END
  END gpio_slow_sel[38]
  PIN gpio_slow_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1278.150 -2.120 1278.430 0.280 ;
    END
  END gpio_slow_sel[39]
  PIN gpio_slow_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 980.115 3168.750 980.465 ;
    END
  END gpio_slow_sel[3]
  PIN gpio_slow_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1552.150 -2.120 1552.430 0.280 ;
    END
  END gpio_slow_sel[40]
  PIN gpio_slow_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1826.150 -2.120 1826.430 0.280 ;
    END
  END gpio_slow_sel[41]
  PIN gpio_slow_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2100.150 -2.120 2100.430 0.280 ;
    END
  END gpio_slow_sel[42]
  PIN gpio_slow_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2374.150 -2.120 2374.430 0.280 ;
    END
  END gpio_slow_sel[43]
  PIN gpio_slow_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1205.115 3168.750 1205.465 ;
    END
  END gpio_slow_sel[4]
  PIN gpio_slow_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1430.115 3168.750 1430.465 ;
    END
  END gpio_slow_sel[5]
  PIN gpio_slow_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1656.115 3168.750 1656.465 ;
    END
  END gpio_slow_sel[6]
  PIN gpio_slow_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2542.115 3168.750 2542.465 ;
    END
  END gpio_slow_sel[7]
  PIN gpio_slow_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2768.115 3168.750 2768.465 ;
    END
  END gpio_slow_sel[8]
  PIN gpio_slow_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2993.115 3168.750 2993.465 ;
    END
  END gpio_slow_sel[9]
  PIN gpio_vtrip_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 358.315 3168.750 358.665 ;
    END
  END gpio_vtrip_sel[0]
  PIN gpio_vtrip_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3274.315 3168.750 3274.665 ;
    END
  END gpio_vtrip_sel[10]
  PIN gpio_vtrip_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3499.315 3168.750 3499.665 ;
    END
  END gpio_vtrip_sel[11]
  PIN gpio_vtrip_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3724.315 3168.750 3724.665 ;
    END
  END gpio_vtrip_sel[12]
  PIN gpio_vtrip_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4170.315 3168.750 4170.665 ;
    END
  END gpio_vtrip_sel[13]
  PIN gpio_vtrip_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 4616.315 3168.750 4616.665 ;
    END
  END gpio_vtrip_sel[14]
  PIN gpio_vtrip_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2930.000 4766.350 2930.280 4768.750 ;
    END
  END gpio_vtrip_sel[15]
  PIN gpio_vtrip_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2421.000 4766.350 2421.280 4768.750 ;
    END
  END gpio_vtrip_sel[16]
  PIN gpio_vtrip_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2164.000 4766.350 2164.280 4768.750 ;
    END
  END gpio_vtrip_sel[17]
  PIN gpio_vtrip_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1719.000 4766.350 1719.280 4768.750 ;
    END
  END gpio_vtrip_sel[18]
  PIN gpio_vtrip_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1210.000 4766.350 1210.280 4768.750 ;
    END
  END gpio_vtrip_sel[19]
  PIN gpio_vtrip_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 584.315 3168.750 584.665 ;
    END
  END gpio_vtrip_sel[1]
  PIN gpio_vtrip_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 952.000 4766.350 952.280 4768.750 ;
    END
  END gpio_vtrip_sel[20]
  PIN gpio_vtrip_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 695.000 4766.350 695.280 4768.750 ;
    END
  END gpio_vtrip_sel[21]
  PIN gpio_vtrip_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 438.000 4766.350 438.280 4768.750 ;
    END
  END gpio_vtrip_sel[22]
  PIN gpio_vtrip_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 181.000 4766.350 181.280 4768.750 ;
    END
  END gpio_vtrip_sel[23]
  PIN gpio_vtrip_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 4570.965 0.280 4571.315 ;
    END
  END gpio_vtrip_sel[24]
  PIN gpio_vtrip_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3721.965 0.280 3722.315 ;
    END
  END gpio_vtrip_sel[25]
  PIN gpio_vtrip_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3505.965 0.280 3506.315 ;
    END
  END gpio_vtrip_sel[26]
  PIN gpio_vtrip_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3289.965 0.280 3290.315 ;
    END
  END gpio_vtrip_sel[27]
  PIN gpio_vtrip_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 3073.965 0.280 3074.315 ;
    END
  END gpio_vtrip_sel[28]
  PIN gpio_vtrip_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2857.965 0.280 2858.315 ;
    END
  END gpio_vtrip_sel[29]
  PIN gpio_vtrip_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 809.315 3168.750 809.665 ;
    END
  END gpio_vtrip_sel[2]
  PIN gpio_vtrip_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2641.965 0.280 2642.315 ;
    END
  END gpio_vtrip_sel[30]
  PIN gpio_vtrip_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 2425.965 0.280 2426.315 ;
    END
  END gpio_vtrip_sel[31]
  PIN gpio_vtrip_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1787.965 0.280 1788.315 ;
    END
  END gpio_vtrip_sel[32]
  PIN gpio_vtrip_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1571.965 0.280 1572.315 ;
    END
  END gpio_vtrip_sel[33]
  PIN gpio_vtrip_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1355.965 0.280 1356.315 ;
    END
  END gpio_vtrip_sel[34]
  PIN gpio_vtrip_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 1139.965 0.280 1140.315 ;
    END
  END gpio_vtrip_sel[35]
  PIN gpio_vtrip_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 923.960 0.280 924.320 ;
    END
  END gpio_vtrip_sel[36]
  PIN gpio_vtrip_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.120 707.960 0.280 708.320 ;
    END
  END gpio_vtrip_sel[37]
  PIN gpio_vtrip_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 790.350 -2.120 790.630 0.280 ;
    END
  END gpio_vtrip_sel[38]
  PIN gpio_vtrip_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1333.350 -2.120 1333.630 0.280 ;
    END
  END gpio_vtrip_sel[39]
  PIN gpio_vtrip_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1035.315 3168.750 1035.665 ;
    END
  END gpio_vtrip_sel[3]
  PIN gpio_vtrip_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1607.350 -2.120 1607.630 0.280 ;
    END
  END gpio_vtrip_sel[40]
  PIN gpio_vtrip_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1881.350 -2.120 1881.630 0.280 ;
    END
  END gpio_vtrip_sel[41]
  PIN gpio_vtrip_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2155.350 -2.120 2155.630 0.280 ;
    END
  END gpio_vtrip_sel[42]
  PIN gpio_vtrip_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2429.350 -2.120 2429.630 0.280 ;
    END
  END gpio_vtrip_sel[43]
  PIN gpio_vtrip_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1260.315 3168.750 1260.665 ;
    END
  END gpio_vtrip_sel[4]
  PIN gpio_vtrip_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1485.315 3168.750 1485.665 ;
    END
  END gpio_vtrip_sel[5]
  PIN gpio_vtrip_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 1711.315 3168.750 1711.665 ;
    END
  END gpio_vtrip_sel[6]
  PIN gpio_vtrip_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2597.315 3168.750 2597.665 ;
    END
  END gpio_vtrip_sel[7]
  PIN gpio_vtrip_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 2823.315 3168.750 2823.665 ;
    END
  END gpio_vtrip_sel[8]
  PIN gpio_vtrip_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3166.350 3048.315 3168.750 3048.665 ;
    END
  END gpio_vtrip_sel[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3025.410 -1.300 3025.670 0.280 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3036.610 -1.300 3036.870 0.280 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3037.730 -1.300 3037.990 0.280 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3038.850 -1.300 3039.110 0.280 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3039.970 -1.300 3040.230 0.280 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3041.090 -1.300 3041.350 0.280 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3042.210 -1.300 3042.470 0.280 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3043.330 -1.300 3043.590 0.280 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3044.450 -1.300 3044.710 0.280 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3045.570 -1.300 3045.830 0.280 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3046.690 -1.300 3046.950 0.280 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3026.530 -1.300 3026.790 0.280 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3047.810 -1.300 3048.070 0.280 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3048.930 -1.300 3049.190 0.280 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3050.050 -1.300 3050.310 0.280 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3051.170 -1.300 3051.430 0.280 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3052.290 -1.300 3052.550 0.280 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3053.410 -1.300 3053.670 0.280 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3054.530 -1.300 3054.790 0.280 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3055.650 -1.300 3055.910 0.280 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3056.770 -1.300 3057.030 0.280 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3057.890 -1.300 3058.150 0.280 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3027.650 -1.300 3027.910 0.280 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3059.010 -1.300 3059.270 0.280 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3060.130 -1.300 3060.390 0.280 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3028.770 -1.300 3029.030 0.280 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3029.890 -1.300 3030.150 0.280 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3031.010 -1.300 3031.270 0.280 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3032.130 -1.300 3032.390 0.280 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3033.250 -1.300 3033.510 0.280 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3034.370 -1.300 3034.630 0.280 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 3035.490 -1.300 3035.750 0.280 ;
    END
  END mask_rev[9]
  PIN por_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.420 266.860 0.280 267.210 ;
    END
  END por_l
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -1.420 265.735 0.280 266.085 ;
    END
  END porb_h
  PIN porb_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT -1.420 267.975 0.280 268.325 ;
    END
  END porb_l
  PIN resetb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.855 -0.450 498.185 0.280 ;
    END
  END resetb_h
  PIN resetb_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 550.820 -0.580 551.100 0.280 ;
    END
  END resetb_l
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.020 24.800 44.020 4740.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 24.020 24.800 3142.620 44.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 24.020 4720.640 3142.620 4740.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 3122.620 24.800 3142.620 4740.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.250 2.400 61.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.250 2.400 101.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.250 2.400 141.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.250 2.400 181.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 215.250 2.400 221.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 255.250 2.400 261.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 295.250 2.400 301.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.250 2.400 341.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 375.250 2.400 381.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 415.250 2.400 421.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 455.250 2.400 461.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.250 2.400 501.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.250 2.400 541.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.250 2.400 581.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.250 3447.990 581.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 615.250 2.400 621.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 615.250 3447.990 621.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.250 2.400 661.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 655.250 3447.990 661.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 695.250 2.400 701.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 695.250 3447.990 701.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 735.250 2.400 741.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 735.250 3447.990 741.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.250 2.400 781.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.250 3447.990 781.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.250 2.400 821.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.250 3447.990 821.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 855.250 2.400 861.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 855.250 3447.990 861.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 895.250 2.400 901.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 895.250 3447.990 901.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 935.250 2.400 941.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 935.250 3447.990 941.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 975.250 2.400 981.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 975.250 3447.990 981.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.250 2.400 1021.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.250 3447.990 1021.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.250 2.400 1061.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.250 3447.990 1061.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.250 2.400 1101.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.250 3447.990 1101.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1135.250 2.400 1141.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1135.250 3447.990 1141.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1175.250 2.400 1181.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1175.250 3447.990 1181.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1215.250 2.400 1221.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1215.250 3447.990 1221.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1255.250 2.400 1261.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1255.250 3447.990 1261.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.250 2.400 1301.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.250 3447.990 1301.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1335.250 2.400 1341.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1335.250 3447.990 1341.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.250 2.400 1381.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.250 3447.990 1381.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1415.250 2.400 1421.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1415.250 3447.990 1421.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1455.250 2.400 1461.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1455.250 3447.990 1461.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1495.250 2.400 1501.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1495.250 3447.990 1501.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1535.250 2.400 1541.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1535.250 3447.990 1541.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.250 2.400 1581.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.250 3447.990 1581.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1615.250 2.400 1621.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1615.250 3447.990 1621.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.250 2.400 1661.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.250 3447.990 1661.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1695.250 2.400 1701.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1695.250 3447.990 1701.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.250 2.400 1741.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.250 3447.990 1741.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1775.250 2.400 1781.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1775.250 3447.990 1781.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1815.250 2.400 1821.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1815.250 3447.990 1821.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1855.250 2.400 1861.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1855.250 3447.990 1861.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1895.250 2.400 1901.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1895.250 3447.990 1901.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.250 2.400 1941.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.250 3447.990 1941.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1975.250 2.400 1981.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1975.250 3447.990 1981.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2015.250 2.400 2021.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2015.250 3447.990 2021.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.250 2.400 2061.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.250 3447.990 2061.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2095.250 2.400 2101.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2095.250 3447.990 2101.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2135.250 2.400 2141.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2135.250 3447.990 2141.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.250 2.400 2181.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.250 3447.990 2181.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.250 2.400 2221.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.250 3447.990 2221.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.250 2.400 2261.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.250 3447.990 2261.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2295.250 2.400 2301.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2295.250 3447.990 2301.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2335.250 2.400 2341.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2335.250 3447.990 2341.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.250 2.400 2381.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.250 3447.990 2381.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2415.250 2.400 2421.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2415.250 3447.990 2421.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2455.250 2.400 2461.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2455.250 3447.990 2461.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2495.250 2.400 2501.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2495.250 3447.990 2501.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2535.250 2.400 2541.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2535.250 3447.990 2541.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2575.250 2.400 2581.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2575.250 3447.990 2581.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2615.250 2.400 2621.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2615.250 3447.990 2621.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2655.250 2.400 2661.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2655.250 3447.990 2661.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2695.250 2.400 2701.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2695.250 3447.990 2701.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2735.250 2.400 2741.650 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2735.250 3447.990 2741.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2775.250 2.400 2781.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2815.250 2.400 2821.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2855.250 2.400 2861.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2895.250 2.400 2901.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2935.250 2.400 2941.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2975.250 2.400 2981.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3015.250 2.400 3021.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3055.250 2.400 3061.650 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3095.250 2.400 3101.650 4763.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 60.430 3165.020 66.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 100.430 3165.020 106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 140.430 3165.020 146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 180.430 3165.020 186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 220.430 3165.020 226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 260.430 3165.020 266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 300.430 3165.020 306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 340.430 3165.020 346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 380.430 3165.020 386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 420.430 3165.020 426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 460.430 3165.020 466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 500.430 3165.020 506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 540.430 3165.020 546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 580.430 3165.020 586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 620.430 3165.020 626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 660.430 3165.020 666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 700.430 3165.020 706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 740.430 3165.020 746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 780.430 3165.020 786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 820.430 3165.020 826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 860.430 3165.020 866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 900.430 3165.020 906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 940.430 3165.020 946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 980.430 3165.020 986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1020.430 3165.020 1026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1060.430 3165.020 1066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1100.430 3165.020 1106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1140.430 3165.020 1146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1180.430 3165.020 1186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1220.430 3165.020 1226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1260.430 3165.020 1266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1300.430 3165.020 1306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1340.430 3165.020 1346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1380.430 3165.020 1386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1420.430 3165.020 1426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1460.430 3165.020 1466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1500.430 3165.020 1506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1540.430 3165.020 1546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1580.430 3165.020 1586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1620.430 3165.020 1626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1660.430 3165.020 1666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1700.430 3165.020 1706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1740.430 3165.020 1746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1780.430 3165.020 1786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1820.430 3165.020 1826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1860.430 3165.020 1866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1900.430 3165.020 1906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1940.430 3165.020 1946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1980.430 3165.020 1986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2020.430 3165.020 2026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2060.430 3165.020 2066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2100.430 3165.020 2106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2140.430 3165.020 2146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2180.430 3165.020 2186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2220.430 3165.020 2226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2260.430 3165.020 2266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2300.430 3165.020 2306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2340.430 3165.020 2346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2380.430 3165.020 2386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2420.430 3165.020 2426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2460.430 3165.020 2466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2500.430 623.860 2506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2540.430 623.860 2546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2580.430 623.860 2586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2620.430 623.860 2626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2660.430 623.860 2666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2700.430 623.860 2706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2740.430 623.860 2746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2780.430 623.860 2786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2820.430 623.860 2826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2860.430 623.860 2866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2900.430 623.860 2906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2940.430 623.860 2946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2980.430 623.860 2986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3020.430 623.860 3026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3060.430 623.860 3066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3100.430 623.860 3106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3140.430 623.860 3146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3180.430 623.860 3186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3220.430 623.860 3226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3260.430 623.860 3266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3300.430 623.860 3306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3340.430 623.860 3346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3380.430 623.860 3386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3420.430 623.860 3426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3460.430 3165.020 3466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3500.430 3165.020 3506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3540.430 3165.020 3546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3580.430 3165.020 3586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3620.430 3165.020 3626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3660.430 3165.020 3666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3700.430 3165.020 3706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3740.430 3165.020 3746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3780.430 3165.020 3786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3820.430 3165.020 3826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3860.430 3165.020 3866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3900.430 3165.020 3906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3940.430 3165.020 3946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3980.430 3165.020 3986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4020.430 3165.020 4026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4060.430 3165.020 4066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4100.430 3165.020 4106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4140.430 3165.020 4146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4180.430 3165.020 4186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4220.430 3165.020 4226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4260.430 3165.020 4266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4300.430 3165.020 4306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4340.430 3165.020 4346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4380.430 3165.020 4386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4420.430 3165.020 4426.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4460.430 3165.020 4466.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4500.430 3165.020 4506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4540.430 3165.020 4546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4580.430 3165.020 4586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4620.430 3165.020 4626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4660.430 3165.020 4666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4700.430 3165.020 4706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2500.430 3165.020 2506.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2540.430 3165.020 2546.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2580.430 3165.020 2586.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2620.430 3165.020 2626.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2660.430 3165.020 2666.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2700.430 3165.020 2706.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2740.430 3165.020 2746.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2780.430 3165.020 2786.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2820.430 3165.020 2826.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2860.430 3165.020 2866.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2900.430 3165.020 2906.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2940.430 3165.020 2946.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2980.430 3165.020 2986.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3020.430 3165.020 3026.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3060.430 3165.020 3066.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3100.430 3165.020 3106.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3140.430 3165.020 3146.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3180.430 3165.020 3186.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3220.430 3165.020 3226.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3260.430 3165.020 3266.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3300.430 3165.020 3306.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3340.430 3165.020 3346.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3380.430 3165.020 3386.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3420.430 3165.020 3426.830 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1.620 2.400 21.620 4763.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2.400 3165.020 22.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4743.040 3165.020 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3145.020 2.400 3165.020 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.850 2.400 71.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.850 2.400 111.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.850 2.400 151.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.850 2.400 191.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.850 2.400 231.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.850 2.400 271.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.850 2.400 311.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.850 2.400 351.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.850 2.400 391.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.850 2.400 431.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.850 2.400 471.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.850 2.400 511.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.850 2.400 551.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 584.850 2.400 591.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 584.850 3447.990 591.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.850 2.400 631.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.850 3447.990 631.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.850 2.400 671.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 664.850 3447.990 671.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.850 2.400 711.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.850 3447.990 711.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.850 2.400 751.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.850 3447.990 751.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.850 2.400 791.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.850 3447.990 791.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 824.850 2.400 831.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 824.850 3447.990 831.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.850 2.400 871.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.850 3447.990 871.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.850 2.400 911.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.850 3447.990 911.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 944.850 2.400 951.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 944.850 3447.990 951.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 984.850 2.400 991.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 984.850 3447.990 991.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.850 2.400 1031.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.850 3447.990 1031.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1064.850 2.400 1071.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1064.850 3447.990 1071.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1104.850 2.400 1111.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1104.850 3447.990 1111.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.850 2.400 1151.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.850 3447.990 1151.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.850 2.400 1191.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.850 3447.990 1191.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.850 2.400 1231.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.850 3447.990 1231.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.850 2.400 1271.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1264.850 3447.990 1271.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.850 2.400 1311.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.850 3447.990 1311.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1344.850 2.400 1351.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1344.850 3447.990 1351.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1384.850 2.400 1391.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1384.850 3447.990 1391.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1424.850 2.400 1431.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1424.850 3447.990 1431.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.850 2.400 1471.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1464.850 3447.990 1471.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.850 2.400 1511.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.850 3447.990 1511.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.850 2.400 1551.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.850 3447.990 1551.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.850 2.400 1591.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.850 3447.990 1591.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1624.850 2.400 1631.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1624.850 3447.990 1631.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.850 2.400 1671.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.850 3447.990 1671.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1704.850 2.400 1711.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1704.850 3447.990 1711.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1744.850 2.400 1751.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1744.850 3447.990 1751.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1784.850 2.400 1791.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1784.850 3447.990 1791.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1824.850 2.400 1831.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1824.850 3447.990 1831.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.850 2.400 1871.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.850 3447.990 1871.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.850 2.400 1911.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.850 3447.990 1911.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1944.850 2.400 1951.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1944.850 3447.990 1951.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.850 2.400 1991.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1984.850 3447.990 1991.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.850 2.400 2031.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.850 3447.990 2031.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2064.850 2.400 2071.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2064.850 3447.990 2071.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2104.850 2.400 2111.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2104.850 3447.990 2111.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.850 2.400 2151.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.850 3447.990 2151.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.850 2.400 2191.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.850 3447.990 2191.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.850 2.400 2231.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.850 3447.990 2231.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2264.850 2.400 2271.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2264.850 3447.990 2271.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.850 2.400 2311.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.850 3447.990 2311.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.850 2.400 2351.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2344.850 3447.990 2351.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2384.850 2.400 2391.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2384.850 3447.990 2391.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.850 2.400 2431.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.850 3447.990 2431.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.850 2.400 2471.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.850 3447.990 2471.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.850 2.400 2511.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.850 3447.990 2511.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2544.850 2.400 2551.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2544.850 3447.990 2551.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.850 2.400 2591.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.850 3447.990 2591.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.850 2.400 2631.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.850 3447.990 2631.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.850 2.400 2671.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2664.850 3447.990 2671.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.850 2.400 2711.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.850 3447.990 2711.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2744.850 2.400 2751.250 2050.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2744.850 3447.990 2751.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2784.850 2.400 2791.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2824.850 2.400 2831.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2864.850 2.400 2871.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2904.850 2.400 2911.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2944.850 2.400 2951.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2984.850 2.400 2991.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3024.850 2.400 3031.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3064.850 2.400 3071.250 4763.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 3104.850 2.400 3111.250 4763.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 70.030 3165.020 76.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 110.030 3165.020 116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 150.030 3165.020 156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 190.030 3165.020 196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 230.030 3165.020 236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 270.030 3165.020 276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 310.030 3165.020 316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 350.030 3165.020 356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 390.030 3165.020 396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 430.030 3165.020 436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 470.030 3165.020 476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 510.030 3165.020 516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 550.030 3165.020 556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 590.030 3165.020 596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 630.030 3165.020 636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 670.030 3165.020 676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 710.030 3165.020 716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 750.030 3165.020 756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 790.030 3165.020 796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 830.030 3165.020 836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 870.030 3165.020 876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 910.030 3165.020 916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 950.030 3165.020 956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 990.030 3165.020 996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1030.030 3165.020 1036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1070.030 3165.020 1076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1110.030 3165.020 1116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1150.030 3165.020 1156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1190.030 3165.020 1196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1230.030 3165.020 1236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1270.030 3165.020 1276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1310.030 3165.020 1316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1350.030 3165.020 1356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1390.030 3165.020 1396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1430.030 3165.020 1436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1470.030 3165.020 1476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1510.030 3165.020 1516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1550.030 3165.020 1556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1590.030 3165.020 1596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1630.030 3165.020 1636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1670.030 3165.020 1676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1710.030 3165.020 1716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1750.030 3165.020 1756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1790.030 3165.020 1796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1830.030 3165.020 1836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1870.030 3165.020 1876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1910.030 3165.020 1916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1950.030 3165.020 1956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 1990.030 3165.020 1996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2030.030 3165.020 2036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2070.030 3165.020 2076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2110.030 3165.020 2116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2150.030 3165.020 2156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2190.030 3165.020 2196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2230.030 3165.020 2236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2270.030 3165.020 2276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2310.030 3165.020 2316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2350.030 3165.020 2356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2390.030 3165.020 2396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2430.030 3165.020 2436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2470.030 3165.020 2476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2510.030 623.860 2516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2550.030 623.860 2556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2590.030 623.860 2596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2630.030 623.860 2636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2670.030 623.860 2676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2710.030 623.860 2716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2750.030 623.860 2756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2790.030 623.860 2796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2830.030 623.860 2836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2870.030 623.860 2876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2910.030 623.860 2916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2950.030 623.860 2956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 2990.030 623.860 2996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3030.030 623.860 3036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3070.030 623.860 3076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3110.030 623.860 3116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3150.030 623.860 3156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3190.030 623.860 3196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3230.030 623.860 3236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3270.030 623.860 3276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3310.030 623.860 3316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3350.030 623.860 3356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3390.030 623.860 3396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3430.030 623.860 3436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3470.030 3165.020 3476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3510.030 3165.020 3516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3550.030 3165.020 3556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3590.030 3165.020 3596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3630.030 3165.020 3636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3670.030 3165.020 3676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3710.030 3165.020 3716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3750.030 3165.020 3756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3790.030 3165.020 3796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3830.030 3165.020 3836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3870.030 3165.020 3876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3910.030 3165.020 3916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3950.030 3165.020 3956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 3990.030 3165.020 3996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4030.030 3165.020 4036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4070.030 3165.020 4076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4110.030 3165.020 4116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4150.030 3165.020 4156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4190.030 3165.020 4196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4230.030 3165.020 4236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4270.030 3165.020 4276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4310.030 3165.020 4316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4350.030 3165.020 4356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4390.030 3165.020 4396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4430.030 3165.020 4436.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4470.030 3165.020 4476.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4510.030 3165.020 4516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4550.030 3165.020 4556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4590.030 3165.020 4596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4630.030 3165.020 4636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4670.030 3165.020 4676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.620 4710.030 3165.020 4716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2510.030 3165.020 2516.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2550.030 3165.020 2556.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2590.030 3165.020 2596.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2630.030 3165.020 2636.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2670.030 3165.020 2676.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2710.030 3165.020 2716.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2750.030 3165.020 2756.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2790.030 3165.020 2796.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2830.030 3165.020 2836.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2870.030 3165.020 2876.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2910.030 3165.020 2916.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2950.030 3165.020 2956.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 2990.030 3165.020 2996.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3030.030 3165.020 3036.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3070.030 3165.020 3076.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3110.030 3165.020 3116.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3150.030 3165.020 3156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3190.030 3165.020 3196.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3230.030 3165.020 3236.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3270.030 3165.020 3276.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3310.030 3165.020 3316.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3350.030 3165.020 3356.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3390.030 3165.020 3396.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2406.300 3430.030 3165.020 3436.430 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 40.020 40.715 3126.620 4724.725 ;
      LAYER met1 ;
        RECT 13.870 13.980 3146.330 4750.100 ;
      LAYER met2 ;
        RECT 13.890 4766.070 137.210 4766.530 ;
        RECT 138.070 4766.070 147.210 4766.530 ;
        RECT 148.070 4766.070 171.520 4766.530 ;
        RECT 172.360 4766.070 174.280 4766.530 ;
        RECT 175.120 4766.070 177.500 4766.530 ;
        RECT 178.340 4766.070 180.720 4766.530 ;
        RECT 181.560 4766.070 189.920 4766.530 ;
        RECT 190.760 4766.070 192.680 4766.530 ;
        RECT 193.520 4766.070 195.900 4766.530 ;
        RECT 196.740 4766.070 199.120 4766.530 ;
        RECT 199.960 4766.070 211.540 4766.530 ;
        RECT 212.380 4766.070 214.300 4766.530 ;
        RECT 215.140 4766.070 217.520 4766.530 ;
        RECT 218.360 4766.070 220.740 4766.530 ;
        RECT 221.580 4766.070 223.500 4766.530 ;
        RECT 224.340 4766.070 226.720 4766.530 ;
        RECT 227.560 4766.070 232.700 4766.530 ;
        RECT 233.540 4766.070 235.920 4766.530 ;
        RECT 236.760 4766.070 245.120 4766.530 ;
        RECT 245.960 4766.070 393.210 4766.530 ;
        RECT 394.070 4766.070 403.210 4766.530 ;
        RECT 404.070 4766.070 428.520 4766.530 ;
        RECT 429.360 4766.070 431.280 4766.530 ;
        RECT 432.120 4766.070 434.500 4766.530 ;
        RECT 435.340 4766.070 437.720 4766.530 ;
        RECT 438.560 4766.070 446.920 4766.530 ;
        RECT 447.760 4766.070 449.680 4766.530 ;
        RECT 450.520 4766.070 452.900 4766.530 ;
        RECT 453.740 4766.070 456.120 4766.530 ;
        RECT 456.960 4766.070 468.540 4766.530 ;
        RECT 469.380 4766.070 471.300 4766.530 ;
        RECT 472.140 4766.070 474.520 4766.530 ;
        RECT 475.360 4766.070 477.740 4766.530 ;
        RECT 478.580 4766.070 480.500 4766.530 ;
        RECT 481.340 4766.070 483.720 4766.530 ;
        RECT 484.560 4766.070 489.700 4766.530 ;
        RECT 490.540 4766.070 492.920 4766.530 ;
        RECT 493.760 4766.070 502.120 4766.530 ;
        RECT 502.960 4766.070 649.210 4766.530 ;
        RECT 650.070 4766.070 659.210 4766.530 ;
        RECT 660.070 4766.070 685.520 4766.530 ;
        RECT 686.360 4766.070 688.280 4766.530 ;
        RECT 689.120 4766.070 691.500 4766.530 ;
        RECT 692.340 4766.070 694.720 4766.530 ;
        RECT 695.560 4766.070 703.920 4766.530 ;
        RECT 704.760 4766.070 706.680 4766.530 ;
        RECT 707.520 4766.070 709.900 4766.530 ;
        RECT 710.740 4766.070 713.120 4766.530 ;
        RECT 713.960 4766.070 725.540 4766.530 ;
        RECT 726.380 4766.070 728.300 4766.530 ;
        RECT 729.140 4766.070 731.520 4766.530 ;
        RECT 732.360 4766.070 734.740 4766.530 ;
        RECT 735.580 4766.070 737.500 4766.530 ;
        RECT 738.340 4766.070 740.720 4766.530 ;
        RECT 741.560 4766.070 746.700 4766.530 ;
        RECT 747.540 4766.070 749.920 4766.530 ;
        RECT 750.760 4766.070 759.120 4766.530 ;
        RECT 759.960 4766.070 905.210 4766.530 ;
        RECT 906.070 4766.070 915.210 4766.530 ;
        RECT 916.070 4766.070 942.520 4766.530 ;
        RECT 943.360 4766.070 945.280 4766.530 ;
        RECT 946.120 4766.070 948.500 4766.530 ;
        RECT 949.340 4766.070 951.720 4766.530 ;
        RECT 952.560 4766.070 960.920 4766.530 ;
        RECT 961.760 4766.070 963.680 4766.530 ;
        RECT 964.520 4766.070 966.900 4766.530 ;
        RECT 967.740 4766.070 970.120 4766.530 ;
        RECT 970.960 4766.070 982.540 4766.530 ;
        RECT 983.380 4766.070 985.300 4766.530 ;
        RECT 986.140 4766.070 988.520 4766.530 ;
        RECT 989.360 4766.070 991.740 4766.530 ;
        RECT 992.580 4766.070 994.500 4766.530 ;
        RECT 995.340 4766.070 997.720 4766.530 ;
        RECT 998.560 4766.070 1003.700 4766.530 ;
        RECT 1004.540 4766.070 1006.920 4766.530 ;
        RECT 1007.760 4766.070 1016.120 4766.530 ;
        RECT 1016.960 4766.070 1161.210 4766.530 ;
        RECT 1162.070 4766.070 1171.210 4766.530 ;
        RECT 1172.070 4766.070 1200.520 4766.530 ;
        RECT 1201.360 4766.070 1203.280 4766.530 ;
        RECT 1204.120 4766.070 1206.500 4766.530 ;
        RECT 1207.340 4766.070 1209.720 4766.530 ;
        RECT 1210.560 4766.070 1218.920 4766.530 ;
        RECT 1219.760 4766.070 1221.680 4766.530 ;
        RECT 1222.520 4766.070 1224.900 4766.530 ;
        RECT 1225.740 4766.070 1228.120 4766.530 ;
        RECT 1228.960 4766.070 1240.540 4766.530 ;
        RECT 1241.380 4766.070 1243.300 4766.530 ;
        RECT 1244.140 4766.070 1246.520 4766.530 ;
        RECT 1247.360 4766.070 1249.740 4766.530 ;
        RECT 1250.580 4766.070 1252.500 4766.530 ;
        RECT 1253.340 4766.070 1255.720 4766.530 ;
        RECT 1256.560 4766.070 1261.700 4766.530 ;
        RECT 1262.540 4766.070 1264.920 4766.530 ;
        RECT 1265.760 4766.070 1274.120 4766.530 ;
        RECT 1274.960 4766.070 1683.210 4766.530 ;
        RECT 1684.070 4766.070 1693.210 4766.530 ;
        RECT 1694.070 4766.070 1709.520 4766.530 ;
        RECT 1710.360 4766.070 1712.280 4766.530 ;
        RECT 1713.120 4766.070 1715.500 4766.530 ;
        RECT 1716.340 4766.070 1718.720 4766.530 ;
        RECT 1719.560 4766.070 1727.920 4766.530 ;
        RECT 1728.760 4766.070 1730.680 4766.530 ;
        RECT 1731.520 4766.070 1733.900 4766.530 ;
        RECT 1734.740 4766.070 1737.120 4766.530 ;
        RECT 1737.960 4766.070 1749.540 4766.530 ;
        RECT 1750.380 4766.070 1752.300 4766.530 ;
        RECT 1753.140 4766.070 1755.520 4766.530 ;
        RECT 1756.360 4766.070 1758.740 4766.530 ;
        RECT 1759.580 4766.070 1761.500 4766.530 ;
        RECT 1762.340 4766.070 1764.720 4766.530 ;
        RECT 1765.560 4766.070 1770.700 4766.530 ;
        RECT 1771.540 4766.070 1773.920 4766.530 ;
        RECT 1774.760 4766.070 1783.120 4766.530 ;
        RECT 1783.960 4766.070 2128.210 4766.530 ;
        RECT 2129.070 4766.070 2138.210 4766.530 ;
        RECT 2139.070 4766.070 2154.520 4766.530 ;
        RECT 2155.360 4766.070 2157.280 4766.530 ;
        RECT 2158.120 4766.070 2160.500 4766.530 ;
        RECT 2161.340 4766.070 2163.720 4766.530 ;
        RECT 2164.560 4766.070 2172.920 4766.530 ;
        RECT 2173.760 4766.070 2175.680 4766.530 ;
        RECT 2176.520 4766.070 2178.900 4766.530 ;
        RECT 2179.740 4766.070 2182.120 4766.530 ;
        RECT 2182.960 4766.070 2194.540 4766.530 ;
        RECT 2195.380 4766.070 2197.300 4766.530 ;
        RECT 2198.140 4766.070 2200.520 4766.530 ;
        RECT 2201.360 4766.070 2203.740 4766.530 ;
        RECT 2204.580 4766.070 2206.500 4766.530 ;
        RECT 2207.340 4766.070 2209.720 4766.530 ;
        RECT 2210.560 4766.070 2215.700 4766.530 ;
        RECT 2216.540 4766.070 2218.920 4766.530 ;
        RECT 2219.760 4766.070 2228.120 4766.530 ;
        RECT 2228.960 4766.070 2384.210 4766.530 ;
        RECT 2385.070 4766.070 2394.210 4766.530 ;
        RECT 2395.070 4766.070 2411.520 4766.530 ;
        RECT 2412.360 4766.070 2414.280 4766.530 ;
        RECT 2415.120 4766.070 2417.500 4766.530 ;
        RECT 2418.340 4766.070 2420.720 4766.530 ;
        RECT 2421.560 4766.070 2429.920 4766.530 ;
        RECT 2430.760 4766.070 2432.680 4766.530 ;
        RECT 2433.520 4766.070 2435.900 4766.530 ;
        RECT 2436.740 4766.070 2439.120 4766.530 ;
        RECT 2439.960 4766.070 2451.540 4766.530 ;
        RECT 2452.380 4766.070 2454.300 4766.530 ;
        RECT 2455.140 4766.070 2457.520 4766.530 ;
        RECT 2458.360 4766.070 2460.740 4766.530 ;
        RECT 2461.580 4766.070 2463.500 4766.530 ;
        RECT 2464.340 4766.070 2466.720 4766.530 ;
        RECT 2467.560 4766.070 2472.700 4766.530 ;
        RECT 2473.540 4766.070 2475.920 4766.530 ;
        RECT 2476.760 4766.070 2485.120 4766.530 ;
        RECT 2485.960 4766.070 2881.210 4766.530 ;
        RECT 2882.070 4766.070 2891.210 4766.530 ;
        RECT 2892.070 4766.070 2920.520 4766.530 ;
        RECT 2921.360 4766.070 2923.280 4766.530 ;
        RECT 2924.120 4766.070 2926.500 4766.530 ;
        RECT 2927.340 4766.070 2929.720 4766.530 ;
        RECT 2930.560 4766.070 2938.920 4766.530 ;
        RECT 2939.760 4766.070 2941.680 4766.530 ;
        RECT 2942.520 4766.070 2944.900 4766.530 ;
        RECT 2945.740 4766.070 2948.120 4766.530 ;
        RECT 2948.960 4766.070 2960.540 4766.530 ;
        RECT 2961.380 4766.070 2963.300 4766.530 ;
        RECT 2964.140 4766.070 2966.520 4766.530 ;
        RECT 2967.360 4766.070 2969.740 4766.530 ;
        RECT 2970.580 4766.070 2972.500 4766.530 ;
        RECT 2973.340 4766.070 2975.720 4766.530 ;
        RECT 2976.560 4766.070 2981.700 4766.530 ;
        RECT 2982.540 4766.070 2984.920 4766.530 ;
        RECT 2985.760 4766.070 2994.120 4766.530 ;
        RECT 2994.960 4766.070 3146.310 4766.530 ;
        RECT 13.890 0.565 3146.310 4766.070 ;
        RECT 13.890 0.560 818.675 0.565 ;
        RECT 13.890 0.070 497.575 0.560 ;
        RECT 498.465 0.070 550.540 0.560 ;
        RECT 551.380 0.070 725.670 0.560 ;
        RECT 726.510 0.070 734.870 0.560 ;
        RECT 735.710 0.070 738.090 0.560 ;
        RECT 738.930 0.070 744.070 0.560 ;
        RECT 744.910 0.070 747.290 0.560 ;
        RECT 748.130 0.070 750.050 0.560 ;
        RECT 750.890 0.070 753.270 0.560 ;
        RECT 754.110 0.070 756.490 0.560 ;
        RECT 757.330 0.070 759.250 0.560 ;
        RECT 760.090 0.070 771.670 0.560 ;
        RECT 772.510 0.070 774.890 0.560 ;
        RECT 775.730 0.070 778.110 0.560 ;
        RECT 778.950 0.070 780.870 0.560 ;
        RECT 781.710 0.070 790.070 0.560 ;
        RECT 790.910 0.070 793.290 0.560 ;
        RECT 794.130 0.070 796.510 0.560 ;
        RECT 797.350 0.070 799.270 0.560 ;
        RECT 800.110 0.070 802.620 0.560 ;
        RECT 803.440 0.070 818.675 0.560 ;
        RECT 819.495 0.560 3146.310 0.565 ;
        RECT 819.495 0.070 1268.670 0.560 ;
        RECT 1269.510 0.070 1277.870 0.560 ;
        RECT 1278.710 0.070 1281.090 0.560 ;
        RECT 1281.930 0.070 1287.070 0.560 ;
        RECT 1287.910 0.070 1290.290 0.560 ;
        RECT 1291.130 0.070 1293.050 0.560 ;
        RECT 1293.890 0.070 1296.270 0.560 ;
        RECT 1297.110 0.070 1299.490 0.560 ;
        RECT 1300.330 0.070 1302.250 0.560 ;
        RECT 1303.090 0.070 1314.670 0.560 ;
        RECT 1315.510 0.070 1317.890 0.560 ;
        RECT 1318.730 0.070 1321.110 0.560 ;
        RECT 1321.950 0.070 1323.870 0.560 ;
        RECT 1324.710 0.070 1333.070 0.560 ;
        RECT 1333.910 0.070 1336.290 0.560 ;
        RECT 1337.130 0.070 1339.510 0.560 ;
        RECT 1340.350 0.070 1342.270 0.560 ;
        RECT 1343.110 0.070 1345.620 0.560 ;
        RECT 1346.440 0.070 1366.520 0.560 ;
        RECT 1367.340 0.070 1542.670 0.560 ;
        RECT 1543.510 0.070 1551.870 0.560 ;
        RECT 1552.710 0.070 1555.090 0.560 ;
        RECT 1555.930 0.070 1561.070 0.560 ;
        RECT 1561.910 0.070 1564.290 0.560 ;
        RECT 1565.130 0.070 1567.050 0.560 ;
        RECT 1567.890 0.070 1570.270 0.560 ;
        RECT 1571.110 0.070 1573.490 0.560 ;
        RECT 1574.330 0.070 1576.250 0.560 ;
        RECT 1577.090 0.070 1588.670 0.560 ;
        RECT 1589.510 0.070 1591.890 0.560 ;
        RECT 1592.730 0.070 1595.110 0.560 ;
        RECT 1595.950 0.070 1597.870 0.560 ;
        RECT 1598.710 0.070 1607.070 0.560 ;
        RECT 1607.910 0.070 1610.290 0.560 ;
        RECT 1611.130 0.070 1613.510 0.560 ;
        RECT 1614.350 0.070 1616.270 0.560 ;
        RECT 1617.110 0.070 1619.620 0.560 ;
        RECT 1620.440 0.450 1816.670 0.560 ;
        RECT 1620.440 0.070 1640.545 0.450 ;
        RECT 1641.365 0.070 1816.670 0.450 ;
        RECT 1817.510 0.070 1825.870 0.560 ;
        RECT 1826.710 0.070 1829.090 0.560 ;
        RECT 1829.930 0.070 1835.070 0.560 ;
        RECT 1835.910 0.070 1838.290 0.560 ;
        RECT 1839.130 0.070 1841.050 0.560 ;
        RECT 1841.890 0.070 1844.270 0.560 ;
        RECT 1845.110 0.070 1847.490 0.560 ;
        RECT 1848.330 0.070 1850.250 0.560 ;
        RECT 1851.090 0.070 1862.670 0.560 ;
        RECT 1863.510 0.070 1865.890 0.560 ;
        RECT 1866.730 0.070 1869.110 0.560 ;
        RECT 1869.950 0.070 1871.870 0.560 ;
        RECT 1872.710 0.070 1881.070 0.560 ;
        RECT 1881.910 0.070 1884.290 0.560 ;
        RECT 1885.130 0.070 1887.510 0.560 ;
        RECT 1888.350 0.070 1890.270 0.560 ;
        RECT 1891.110 0.070 1893.620 0.560 ;
        RECT 1894.440 0.070 1914.610 0.560 ;
        RECT 1915.430 0.070 2090.670 0.560 ;
        RECT 2091.510 0.070 2099.870 0.560 ;
        RECT 2100.710 0.070 2103.090 0.560 ;
        RECT 2103.930 0.070 2109.070 0.560 ;
        RECT 2109.910 0.070 2112.290 0.560 ;
        RECT 2113.130 0.070 2115.050 0.560 ;
        RECT 2115.890 0.070 2118.270 0.560 ;
        RECT 2119.110 0.070 2121.490 0.560 ;
        RECT 2122.330 0.070 2124.250 0.560 ;
        RECT 2125.090 0.070 2136.670 0.560 ;
        RECT 2137.510 0.070 2139.890 0.560 ;
        RECT 2140.730 0.070 2143.110 0.560 ;
        RECT 2143.950 0.070 2145.870 0.560 ;
        RECT 2146.710 0.070 2155.070 0.560 ;
        RECT 2155.910 0.070 2158.290 0.560 ;
        RECT 2159.130 0.070 2161.510 0.560 ;
        RECT 2162.350 0.070 2164.270 0.560 ;
        RECT 2165.110 0.070 2167.620 0.560 ;
        RECT 2168.440 0.070 2188.610 0.560 ;
        RECT 2189.430 0.070 2364.670 0.560 ;
        RECT 2365.510 0.070 2373.870 0.560 ;
        RECT 2374.710 0.070 2377.090 0.560 ;
        RECT 2377.930 0.070 2383.070 0.560 ;
        RECT 2383.910 0.070 2386.290 0.560 ;
        RECT 2387.130 0.070 2389.050 0.560 ;
        RECT 2389.890 0.070 2392.270 0.560 ;
        RECT 2393.110 0.070 2395.490 0.560 ;
        RECT 2396.330 0.070 2398.250 0.560 ;
        RECT 2399.090 0.070 2410.670 0.560 ;
        RECT 2411.510 0.070 2413.890 0.560 ;
        RECT 2414.730 0.070 2417.110 0.560 ;
        RECT 2417.950 0.070 2419.870 0.560 ;
        RECT 2420.710 0.070 2429.070 0.560 ;
        RECT 2429.910 0.070 2432.290 0.560 ;
        RECT 2433.130 0.070 2435.510 0.560 ;
        RECT 2436.350 0.070 2438.270 0.560 ;
        RECT 2439.110 0.070 2441.620 0.560 ;
        RECT 2442.440 0.070 2462.895 0.560 ;
        RECT 2463.715 0.070 3025.130 0.560 ;
        RECT 3025.950 0.070 3026.250 0.560 ;
        RECT 3027.070 0.070 3027.370 0.560 ;
        RECT 3028.190 0.070 3028.490 0.560 ;
        RECT 3029.310 0.070 3029.610 0.560 ;
        RECT 3030.430 0.070 3030.730 0.560 ;
        RECT 3031.550 0.070 3031.850 0.560 ;
        RECT 3032.670 0.070 3032.970 0.560 ;
        RECT 3033.790 0.070 3034.090 0.560 ;
        RECT 3034.910 0.070 3035.210 0.560 ;
        RECT 3036.030 0.070 3036.330 0.560 ;
        RECT 3037.150 0.070 3037.450 0.560 ;
        RECT 3038.270 0.070 3038.570 0.560 ;
        RECT 3039.390 0.070 3039.690 0.560 ;
        RECT 3040.510 0.070 3040.810 0.560 ;
        RECT 3041.630 0.070 3041.930 0.560 ;
        RECT 3042.750 0.070 3043.050 0.560 ;
        RECT 3043.870 0.070 3044.170 0.560 ;
        RECT 3044.990 0.070 3045.290 0.560 ;
        RECT 3046.110 0.070 3046.410 0.560 ;
        RECT 3047.230 0.070 3047.530 0.560 ;
        RECT 3048.350 0.070 3048.650 0.560 ;
        RECT 3049.470 0.070 3049.770 0.560 ;
        RECT 3050.590 0.070 3050.890 0.560 ;
        RECT 3051.710 0.070 3052.010 0.560 ;
        RECT 3052.830 0.070 3053.130 0.560 ;
        RECT 3053.950 0.070 3054.250 0.560 ;
        RECT 3055.070 0.070 3055.370 0.560 ;
        RECT 3056.190 0.070 3056.490 0.560 ;
        RECT 3057.310 0.070 3057.610 0.560 ;
        RECT 3058.430 0.070 3058.730 0.560 ;
        RECT 3059.550 0.070 3059.850 0.560 ;
        RECT 3060.670 0.070 3146.310 0.560 ;
      LAYER met3 ;
        RECT 0.000 4645.745 3166.630 4724.805 ;
        RECT 0.000 4644.635 3165.950 4645.745 ;
        RECT 0.000 4636.115 3166.630 4644.635 ;
        RECT 0.680 4635.735 3166.630 4636.115 ;
        RECT 0.680 4634.965 3165.950 4635.735 ;
        RECT 0.000 4634.625 3165.950 4634.965 ;
        RECT 0.000 4626.915 3166.630 4634.625 ;
        RECT 0.680 4626.265 3166.630 4626.915 ;
        RECT 0.680 4625.765 3165.950 4626.265 ;
        RECT 0.000 4625.115 3165.950 4625.765 ;
        RECT 0.000 4623.695 3166.630 4625.115 ;
        RECT 0.680 4623.505 3166.630 4623.695 ;
        RECT 0.680 4622.545 3165.950 4623.505 ;
        RECT 0.000 4622.355 3165.950 4622.545 ;
        RECT 0.000 4620.285 3166.630 4622.355 ;
        RECT 0.000 4619.135 3165.950 4620.285 ;
        RECT 0.000 4617.715 3166.630 4619.135 ;
        RECT 0.680 4617.065 3166.630 4617.715 ;
        RECT 0.680 4616.565 3165.950 4617.065 ;
        RECT 0.000 4615.915 3165.950 4616.565 ;
        RECT 0.000 4614.495 3166.630 4615.915 ;
        RECT 0.680 4613.345 3166.630 4614.495 ;
        RECT 0.000 4611.735 3166.630 4613.345 ;
        RECT 0.680 4610.585 3166.630 4611.735 ;
        RECT 0.000 4608.515 3166.630 4610.585 ;
        RECT 0.680 4607.865 3166.630 4608.515 ;
        RECT 0.680 4607.365 3165.950 4607.865 ;
        RECT 0.000 4606.715 3165.950 4607.365 ;
        RECT 0.000 4605.295 3166.630 4606.715 ;
        RECT 0.680 4605.105 3166.630 4605.295 ;
        RECT 0.680 4604.145 3165.950 4605.105 ;
        RECT 0.000 4603.955 3165.950 4604.145 ;
        RECT 0.000 4602.535 3166.630 4603.955 ;
        RECT 0.680 4601.885 3166.630 4602.535 ;
        RECT 0.680 4601.385 3165.950 4601.885 ;
        RECT 0.000 4600.735 3165.950 4601.385 ;
        RECT 0.000 4598.665 3166.630 4600.735 ;
        RECT 0.000 4597.515 3165.950 4598.665 ;
        RECT 0.000 4590.115 3166.630 4597.515 ;
        RECT 0.680 4588.965 3166.630 4590.115 ;
        RECT 0.000 4586.895 3166.630 4588.965 ;
        RECT 0.680 4586.245 3166.630 4586.895 ;
        RECT 0.680 4585.745 3165.950 4586.245 ;
        RECT 0.000 4585.095 3165.950 4585.745 ;
        RECT 0.000 4585.050 3166.630 4585.095 ;
        RECT 0.000 4583.675 3166.640 4585.050 ;
        RECT 0.680 4583.390 3166.640 4583.675 ;
        RECT 0.680 4582.525 3165.950 4583.390 ;
        RECT 0.000 4582.335 3165.950 4582.525 ;
        RECT 0.000 4580.915 3166.630 4582.335 ;
        RECT 0.680 4580.265 3166.630 4580.915 ;
        RECT -0.010 4579.990 0.610 4580.165 ;
        RECT -0.010 4579.765 0.290 4579.990 ;
        RECT 0.680 4579.765 3165.950 4580.265 ;
        RECT -0.010 4579.310 3165.950 4579.765 ;
        RECT 0.000 4579.115 3165.950 4579.310 ;
        RECT 0.000 4577.045 3166.630 4579.115 ;
        RECT 0.000 4575.895 3165.950 4577.045 ;
        RECT 0.000 4574.285 3166.630 4575.895 ;
        RECT 0.000 4573.135 3165.950 4574.285 ;
        RECT 0.000 4571.715 3166.630 4573.135 ;
        RECT 0.680 4571.065 3166.630 4571.715 ;
        RECT 0.680 4570.565 3165.950 4571.065 ;
        RECT 0.000 4569.915 3165.950 4570.565 ;
        RECT 0.000 4568.495 3166.630 4569.915 ;
        RECT 0.680 4567.345 3166.630 4568.495 ;
        RECT 0.000 4565.275 3166.630 4567.345 ;
        RECT 0.680 4565.085 3166.630 4565.275 ;
        RECT 0.680 4564.125 3165.950 4565.085 ;
        RECT 0.000 4563.935 3165.950 4564.125 ;
        RECT 0.000 4562.515 3166.630 4563.935 ;
        RECT 0.680 4561.865 3166.630 4562.515 ;
        RECT 0.680 4561.365 3165.950 4561.865 ;
        RECT 0.000 4560.715 3165.950 4561.365 ;
        RECT 0.000 4552.665 3166.630 4560.715 ;
        RECT 0.000 4551.515 3165.950 4552.665 ;
        RECT 0.000 4533.920 3166.630 4551.515 ;
        RECT 0.680 4532.820 3166.630 4533.920 ;
        RECT 0.000 4523.920 3166.630 4532.820 ;
        RECT 0.680 4522.820 3166.630 4523.920 ;
        RECT 0.000 4401.815 3166.630 4522.820 ;
        RECT 0.000 4327.615 3122.620 4401.815 ;
      LAYER met3 ;
        RECT 3122.620 4327.615 3167.855 4401.815 ;
      LAYER met3 ;
        RECT 0.000 4195.745 3166.630 4327.615 ;
        RECT 0.000 4194.635 3165.950 4195.745 ;
        RECT 0.000 4185.735 3166.630 4194.635 ;
        RECT 0.000 4184.625 3165.950 4185.735 ;
        RECT 0.000 4180.265 3166.630 4184.625 ;
        RECT 0.000 4179.115 3165.950 4180.265 ;
        RECT 0.000 4177.505 3166.630 4179.115 ;
        RECT 0.000 4176.355 3165.950 4177.505 ;
        RECT 0.000 4174.285 3166.630 4176.355 ;
        RECT 0.000 4173.135 3165.950 4174.285 ;
        RECT 0.000 4172.290 3166.630 4173.135 ;
        RECT 0.000 4171.065 3166.640 4172.290 ;
        RECT 0.000 4169.915 3165.950 4171.065 ;
        RECT 3166.340 4170.930 3166.640 4171.065 ;
        RECT 3166.030 4170.665 3166.640 4170.930 ;
        RECT 0.000 4161.865 3166.630 4169.915 ;
        RECT 0.000 4160.715 3165.950 4161.865 ;
        RECT 0.000 4159.105 3166.630 4160.715 ;
        RECT 0.000 4157.955 3165.950 4159.105 ;
        RECT 0.000 4155.885 3166.630 4157.955 ;
        RECT 0.000 4154.735 3165.950 4155.885 ;
        RECT 0.000 4152.665 3166.630 4154.735 ;
        RECT 0.000 4151.515 3165.950 4152.665 ;
        RECT 0.000 4140.245 3166.630 4151.515 ;
        RECT 0.000 4139.095 3165.950 4140.245 ;
        RECT 0.000 4137.485 3166.630 4139.095 ;
        RECT 0.000 4136.335 3165.950 4137.485 ;
        RECT 0.000 4134.265 3166.630 4136.335 ;
        RECT 0.000 4133.115 3165.950 4134.265 ;
        RECT 0.000 4131.490 3166.630 4133.115 ;
        RECT 0.000 4131.045 3166.640 4131.490 ;
        RECT 0.000 4129.895 3165.950 4131.045 ;
        RECT 3166.340 4130.810 3166.640 4131.045 ;
        RECT 3166.030 4130.645 3166.640 4130.810 ;
        RECT 0.000 4128.285 3166.630 4129.895 ;
        RECT 0.000 4127.135 3165.950 4128.285 ;
        RECT 0.000 4125.065 3166.630 4127.135 ;
        RECT 0.000 4123.915 3165.950 4125.065 ;
        RECT 0.000 4119.085 3166.630 4123.915 ;
        RECT 0.000 4117.935 3165.950 4119.085 ;
        RECT 0.000 4115.865 3166.630 4117.935 ;
        RECT 0.000 4114.715 3165.950 4115.865 ;
        RECT 3166.030 4114.870 3166.640 4115.115 ;
        RECT 3166.340 4114.715 3166.640 4114.870 ;
        RECT 0.000 4114.190 3166.640 4114.715 ;
        RECT 0.000 4106.665 3166.630 4114.190 ;
        RECT 0.000 4105.515 3165.950 4106.665 ;
        RECT 0.000 3787.115 3166.630 4105.515 ;
        RECT 0.680 3785.965 3166.630 3787.115 ;
        RECT 0.000 3777.915 3166.630 3785.965 ;
        RECT 0.680 3776.765 3166.630 3777.915 ;
        RECT 0.000 3774.695 3166.630 3776.765 ;
        RECT 0.680 3773.545 3166.630 3774.695 ;
        RECT 0.000 3768.715 3166.630 3773.545 ;
        RECT 0.680 3767.565 3166.630 3768.715 ;
        RECT 0.000 3765.495 3166.630 3767.565 ;
        RECT 0.680 3764.345 3166.630 3765.495 ;
        RECT 0.000 3762.735 3166.630 3764.345 ;
        RECT 0.680 3761.585 3166.630 3762.735 ;
        RECT 0.000 3759.515 3166.630 3761.585 ;
        RECT 0.680 3758.365 3166.630 3759.515 ;
        RECT 0.000 3756.295 3166.630 3758.365 ;
        RECT 0.680 3755.145 3166.630 3756.295 ;
        RECT 0.000 3753.535 3166.630 3755.145 ;
        RECT 0.680 3752.385 3166.630 3753.535 ;
        RECT 0.000 3750.745 3166.630 3752.385 ;
        RECT 0.000 3749.635 3165.950 3750.745 ;
        RECT 0.000 3741.170 3166.630 3749.635 ;
        RECT 0.000 3741.115 3166.640 3741.170 ;
        RECT 0.680 3740.735 3166.640 3741.115 ;
        RECT 0.680 3739.965 3165.950 3740.735 ;
        RECT 3166.340 3740.490 3166.640 3740.735 ;
        RECT 3166.030 3740.335 3166.640 3740.490 ;
        RECT 0.000 3739.625 3165.950 3739.965 ;
        RECT 0.000 3737.895 3166.630 3739.625 ;
        RECT 0.680 3736.745 3166.630 3737.895 ;
        RECT 0.000 3734.675 3166.630 3736.745 ;
        RECT 0.680 3734.265 3166.630 3734.675 ;
        RECT 0.680 3733.525 3165.950 3734.265 ;
        RECT 0.000 3733.115 3165.950 3733.525 ;
        RECT 0.000 3731.915 3166.630 3733.115 ;
        RECT 0.680 3731.505 3166.630 3731.915 ;
        RECT 0.680 3730.765 3165.950 3731.505 ;
        RECT 0.000 3730.355 3165.950 3730.765 ;
        RECT 0.000 3728.285 3166.630 3730.355 ;
        RECT 0.000 3727.135 3165.950 3728.285 ;
        RECT 0.000 3725.530 3166.630 3727.135 ;
        RECT 0.000 3725.065 3166.640 3725.530 ;
        RECT 0.000 3723.915 3165.950 3725.065 ;
        RECT 3166.340 3724.850 3166.640 3725.065 ;
        RECT 3166.030 3724.665 3166.640 3724.850 ;
        RECT 0.000 3722.715 3166.630 3723.915 ;
        RECT 0.680 3721.565 3166.630 3722.715 ;
        RECT 0.000 3719.495 3166.630 3721.565 ;
        RECT 0.680 3718.345 3166.630 3719.495 ;
        RECT 0.000 3716.275 3166.630 3718.345 ;
        RECT 0.680 3715.865 3166.630 3716.275 ;
        RECT 0.680 3715.125 3165.950 3715.865 ;
        RECT 0.000 3714.715 3165.950 3715.125 ;
        RECT 0.000 3713.515 3166.630 3714.715 ;
        RECT 0.680 3713.105 3166.630 3713.515 ;
        RECT 0.680 3712.365 3165.950 3713.105 ;
        RECT 0.000 3711.955 3165.950 3712.365 ;
        RECT 0.000 3709.885 3166.630 3711.955 ;
        RECT 0.000 3708.735 3165.950 3709.885 ;
        RECT 0.000 3706.665 3166.630 3708.735 ;
        RECT 0.000 3705.515 3165.950 3706.665 ;
        RECT 0.000 3694.245 3166.630 3705.515 ;
        RECT 0.000 3693.095 3165.950 3694.245 ;
        RECT 0.000 3691.485 3166.630 3693.095 ;
        RECT 0.000 3690.335 3165.950 3691.485 ;
        RECT 3166.030 3690.550 3166.640 3690.735 ;
        RECT 3166.340 3690.335 3166.640 3690.550 ;
        RECT 0.000 3689.870 3166.640 3690.335 ;
        RECT 0.000 3688.810 3166.630 3689.870 ;
        RECT 0.000 3688.265 3166.640 3688.810 ;
        RECT 0.000 3687.115 3165.950 3688.265 ;
        RECT 3166.340 3688.130 3166.640 3688.265 ;
        RECT 3166.030 3687.865 3166.640 3688.130 ;
        RECT 0.000 3685.045 3166.630 3687.115 ;
        RECT 0.000 3683.920 3165.950 3685.045 ;
        RECT 0.680 3683.895 3165.950 3683.920 ;
        RECT 0.680 3682.820 3166.630 3683.895 ;
        RECT 0.000 3682.285 3166.630 3682.820 ;
        RECT 0.000 3681.135 3165.950 3682.285 ;
        RECT 0.000 3679.065 3166.630 3681.135 ;
        RECT 0.000 3677.915 3165.950 3679.065 ;
        RECT 0.000 3673.920 3166.630 3677.915 ;
        RECT 0.680 3673.085 3166.630 3673.920 ;
        RECT 0.680 3672.820 3165.950 3673.085 ;
        RECT 0.000 3671.935 3165.950 3672.820 ;
        RECT 0.000 3669.865 3166.630 3671.935 ;
        RECT 0.000 3668.715 3165.950 3669.865 ;
        RECT 0.000 3661.610 3166.630 3668.715 ;
        RECT 0.000 3660.665 3166.640 3661.610 ;
        RECT 0.000 3659.515 3165.950 3660.665 ;
        RECT 3166.340 3660.420 3166.640 3660.665 ;
        RECT 3166.030 3660.265 3166.640 3660.420 ;
        RECT 0.000 3571.115 3166.630 3659.515 ;
        RECT 0.680 3569.965 3166.630 3571.115 ;
        RECT 0.000 3561.915 3166.630 3569.965 ;
        RECT 0.680 3560.765 3166.630 3561.915 ;
        RECT 0.000 3558.695 3166.630 3560.765 ;
        RECT 0.680 3557.545 3166.630 3558.695 ;
        RECT 0.000 3552.715 3166.630 3557.545 ;
        RECT 0.680 3551.565 3166.630 3552.715 ;
        RECT 0.000 3549.495 3166.630 3551.565 ;
        RECT 0.680 3548.345 3166.630 3549.495 ;
        RECT 0.000 3546.735 3166.630 3548.345 ;
        RECT 0.680 3545.585 3166.630 3546.735 ;
        RECT 0.000 3543.970 3166.630 3545.585 ;
        RECT -0.010 3543.515 3166.630 3543.970 ;
        RECT -0.010 3543.290 0.290 3543.515 ;
        RECT -0.010 3543.115 0.610 3543.290 ;
        RECT 0.680 3542.365 3166.630 3543.515 ;
        RECT 0.000 3540.295 3166.630 3542.365 ;
        RECT 0.680 3539.145 3166.630 3540.295 ;
        RECT 0.000 3537.535 3166.630 3539.145 ;
        RECT 0.680 3536.385 3166.630 3537.535 ;
        RECT 0.000 3525.745 3166.630 3536.385 ;
        RECT 0.000 3525.610 3165.950 3525.745 ;
        RECT -0.010 3525.115 3165.950 3525.610 ;
        RECT -0.010 3524.930 0.290 3525.115 ;
        RECT -0.010 3524.715 0.610 3524.930 ;
        RECT 0.680 3524.635 3165.950 3525.115 ;
        RECT 0.680 3523.965 3166.630 3524.635 ;
        RECT 0.000 3521.895 3166.630 3523.965 ;
        RECT 0.680 3520.745 3166.630 3521.895 ;
        RECT 0.000 3518.675 3166.630 3520.745 ;
        RECT 0.680 3517.525 3166.630 3518.675 ;
        RECT 0.000 3515.915 3166.630 3517.525 ;
        RECT 0.680 3515.735 3166.630 3515.915 ;
        RECT 0.680 3514.765 3165.950 3515.735 ;
        RECT 0.000 3514.625 3165.950 3514.765 ;
        RECT 0.000 3509.265 3166.630 3514.625 ;
        RECT 0.000 3508.115 3165.950 3509.265 ;
        RECT 0.000 3506.715 3166.630 3508.115 ;
        RECT 0.680 3506.505 3166.630 3506.715 ;
        RECT 0.680 3505.565 3165.950 3506.505 ;
        RECT 0.000 3505.355 3165.950 3505.565 ;
        RECT 0.000 3503.495 3166.630 3505.355 ;
        RECT 0.680 3503.285 3166.630 3503.495 ;
        RECT 0.680 3502.345 3165.950 3503.285 ;
        RECT 0.000 3502.135 3165.950 3502.345 ;
        RECT 0.000 3500.275 3166.630 3502.135 ;
        RECT 0.680 3500.065 3166.630 3500.275 ;
        RECT 0.680 3499.125 3165.950 3500.065 ;
        RECT 0.000 3498.915 3165.950 3499.125 ;
        RECT 0.000 3497.515 3166.630 3498.915 ;
        RECT 0.680 3496.365 3166.630 3497.515 ;
        RECT 0.000 3490.865 3166.630 3496.365 ;
        RECT 0.000 3489.715 3165.950 3490.865 ;
        RECT 0.000 3488.105 3166.630 3489.715 ;
        RECT 0.000 3486.955 3165.950 3488.105 ;
        RECT 0.000 3484.885 3166.630 3486.955 ;
        RECT 0.000 3483.735 3165.950 3484.885 ;
        RECT 0.000 3481.665 3166.630 3483.735 ;
        RECT 0.000 3480.515 3165.950 3481.665 ;
        RECT 0.000 3469.245 3166.630 3480.515 ;
        RECT 0.000 3468.920 3165.950 3469.245 ;
        RECT 0.680 3468.095 3165.950 3468.920 ;
        RECT 0.680 3467.820 3166.630 3468.095 ;
        RECT 0.000 3466.485 3166.630 3467.820 ;
        RECT 0.000 3465.335 3165.950 3466.485 ;
        RECT 0.000 3463.730 3166.630 3465.335 ;
        RECT 0.000 3463.265 3166.640 3463.730 ;
        RECT 0.000 3462.115 3165.950 3463.265 ;
        RECT 3166.340 3463.050 3166.640 3463.265 ;
        RECT 3166.030 3462.865 3166.640 3463.050 ;
        RECT 0.000 3460.045 3166.630 3462.115 ;
        RECT 0.000 3458.920 3165.950 3460.045 ;
        RECT 0.680 3458.895 3165.950 3458.920 ;
        RECT 0.680 3457.820 3166.630 3458.895 ;
        RECT 0.000 3457.285 3166.630 3457.820 ;
        RECT 0.000 3456.135 3165.950 3457.285 ;
        RECT 0.000 3454.065 3166.630 3456.135 ;
        RECT 0.000 3452.915 3165.950 3454.065 ;
        RECT 0.000 3448.085 3166.630 3452.915 ;
        RECT 0.000 3446.935 3165.950 3448.085 ;
        RECT 0.000 3444.865 3166.630 3446.935 ;
        RECT 0.000 3443.715 3165.950 3444.865 ;
        RECT 0.000 3435.665 3166.630 3443.715 ;
        RECT 0.000 3434.515 3165.950 3435.665 ;
        RECT 0.000 3355.115 3166.630 3434.515 ;
        RECT 0.680 3353.965 3166.630 3355.115 ;
        RECT 0.000 3345.915 3166.630 3353.965 ;
        RECT 0.680 3344.765 3166.630 3345.915 ;
        RECT 0.000 3342.695 3166.630 3344.765 ;
        RECT 0.680 3341.545 3166.630 3342.695 ;
        RECT 0.000 3337.250 3166.630 3341.545 ;
        RECT -0.010 3336.715 3166.630 3337.250 ;
        RECT -0.010 3336.570 0.290 3336.715 ;
        RECT -0.010 3336.315 0.610 3336.570 ;
        RECT 0.680 3335.565 3166.630 3336.715 ;
        RECT 0.000 3333.495 3166.630 3335.565 ;
        RECT 0.680 3332.345 3166.630 3333.495 ;
        RECT 0.000 3330.735 3166.630 3332.345 ;
        RECT 0.680 3329.585 3166.630 3330.735 ;
        RECT 0.000 3327.515 3166.630 3329.585 ;
        RECT 0.680 3326.365 3166.630 3327.515 ;
        RECT 0.000 3324.295 3166.630 3326.365 ;
        RECT 0.680 3323.145 3166.630 3324.295 ;
        RECT 0.000 3321.535 3166.630 3323.145 ;
        RECT -0.010 3320.630 0.610 3320.785 ;
        RECT -0.010 3320.385 0.290 3320.630 ;
        RECT 0.680 3320.385 3166.630 3321.535 ;
        RECT -0.010 3319.950 3166.630 3320.385 ;
        RECT 0.000 3309.115 3166.630 3319.950 ;
        RECT 0.680 3307.965 3166.630 3309.115 ;
        RECT 0.000 3305.895 3166.630 3307.965 ;
        RECT 0.680 3304.745 3166.630 3305.895 ;
        RECT 0.000 3302.675 3166.630 3304.745 ;
        RECT 0.680 3301.525 3166.630 3302.675 ;
        RECT 0.000 3300.745 3166.630 3301.525 ;
        RECT 0.000 3299.915 3165.950 3300.745 ;
        RECT 0.680 3299.635 3165.950 3299.915 ;
        RECT 0.680 3298.765 3166.630 3299.635 ;
        RECT 0.000 3290.735 3166.630 3298.765 ;
        RECT 0.000 3290.715 3165.950 3290.735 ;
        RECT 0.680 3289.625 3165.950 3290.715 ;
        RECT 0.680 3289.565 3166.630 3289.625 ;
        RECT 0.000 3287.495 3166.630 3289.565 ;
        RECT 0.680 3286.345 3166.630 3287.495 ;
        RECT 0.000 3284.275 3166.630 3286.345 ;
        RECT 0.680 3284.265 3166.630 3284.275 ;
        RECT 0.680 3283.125 3165.950 3284.265 ;
        RECT 0.000 3283.115 3165.950 3283.125 ;
        RECT 0.000 3281.515 3166.630 3283.115 ;
        RECT 0.680 3281.505 3166.630 3281.515 ;
        RECT 0.680 3280.365 3165.950 3281.505 ;
        RECT 0.000 3280.355 3165.950 3280.365 ;
        RECT 0.000 3278.285 3166.630 3280.355 ;
        RECT 0.000 3277.135 3165.950 3278.285 ;
        RECT 0.000 3275.065 3166.630 3277.135 ;
        RECT 0.000 3273.915 3165.950 3275.065 ;
        RECT 0.000 3265.865 3166.630 3273.915 ;
        RECT 0.000 3264.715 3165.950 3265.865 ;
        RECT 0.000 3263.105 3166.630 3264.715 ;
        RECT 0.000 3261.955 3165.950 3263.105 ;
        RECT 0.000 3261.090 3166.630 3261.955 ;
        RECT 0.000 3259.885 3166.640 3261.090 ;
        RECT 0.000 3258.735 3165.950 3259.885 ;
        RECT 3166.340 3259.730 3166.640 3259.885 ;
        RECT 3166.030 3259.485 3166.640 3259.730 ;
        RECT 0.000 3256.665 3166.630 3258.735 ;
        RECT 0.000 3255.515 3165.950 3256.665 ;
        RECT 0.000 3253.920 3166.630 3255.515 ;
        RECT 0.680 3252.820 3166.630 3253.920 ;
        RECT 0.000 3247.490 3166.630 3252.820 ;
        RECT 0.000 3244.245 3166.640 3247.490 ;
        RECT 0.000 3243.920 3165.950 3244.245 ;
        RECT 3166.340 3244.090 3166.640 3244.245 ;
        RECT 0.680 3243.095 3165.950 3243.920 ;
        RECT 3166.030 3243.845 3166.640 3244.090 ;
        RECT 0.680 3242.820 3166.630 3243.095 ;
        RECT 0.000 3241.485 3166.630 3242.820 ;
        RECT 0.000 3240.335 3165.950 3241.485 ;
        RECT 0.000 3238.265 3166.630 3240.335 ;
        RECT 0.000 3237.115 3165.950 3238.265 ;
        RECT 0.000 3235.045 3166.630 3237.115 ;
        RECT 0.000 3233.895 3165.950 3235.045 ;
        RECT 0.000 3232.285 3166.630 3233.895 ;
        RECT 0.000 3231.135 3165.950 3232.285 ;
        RECT 0.000 3229.065 3166.630 3231.135 ;
        RECT 0.000 3227.915 3165.950 3229.065 ;
        RECT 3166.030 3228.150 3166.640 3228.315 ;
        RECT 3166.340 3227.915 3166.640 3228.150 ;
        RECT 0.000 3227.470 3166.640 3227.915 ;
        RECT 0.000 3223.085 3166.630 3227.470 ;
        RECT 0.000 3221.935 3165.950 3223.085 ;
        RECT 0.000 3219.865 3166.630 3221.935 ;
        RECT 0.000 3218.715 3165.950 3219.865 ;
        RECT 0.000 3210.665 3166.630 3218.715 ;
        RECT 0.000 3209.515 3165.950 3210.665 ;
        RECT 0.000 3139.115 3166.630 3209.515 ;
        RECT 0.680 3137.965 3166.630 3139.115 ;
        RECT 0.000 3129.915 3166.630 3137.965 ;
        RECT 0.680 3128.765 3166.630 3129.915 ;
        RECT 0.000 3126.695 3166.630 3128.765 ;
        RECT 0.680 3125.545 3166.630 3126.695 ;
        RECT 0.000 3120.715 3166.630 3125.545 ;
        RECT 0.680 3119.565 3166.630 3120.715 ;
        RECT 0.000 3117.495 3166.630 3119.565 ;
        RECT 0.680 3116.345 3166.630 3117.495 ;
        RECT 0.000 3114.735 3166.630 3116.345 ;
        RECT 0.680 3113.585 3166.630 3114.735 ;
        RECT 0.000 3111.515 3166.630 3113.585 ;
        RECT 0.680 3110.365 3166.630 3111.515 ;
        RECT 0.000 3108.770 3166.630 3110.365 ;
        RECT -0.010 3108.295 3166.630 3108.770 ;
        RECT -0.010 3108.090 0.290 3108.295 ;
        RECT -0.010 3107.895 0.610 3108.090 ;
        RECT 0.680 3107.145 3166.630 3108.295 ;
        RECT 0.000 3105.535 3166.630 3107.145 ;
        RECT 0.680 3104.385 3166.630 3105.535 ;
        RECT 0.000 3093.115 3166.630 3104.385 ;
        RECT 0.680 3091.965 3166.630 3093.115 ;
        RECT 0.000 3089.895 3166.630 3091.965 ;
        RECT 0.680 3088.745 3166.630 3089.895 ;
        RECT 0.000 3086.675 3166.630 3088.745 ;
        RECT 0.680 3085.525 3166.630 3086.675 ;
        RECT 0.000 3083.915 3166.630 3085.525 ;
        RECT 0.680 3082.765 3166.630 3083.915 ;
        RECT 0.000 3075.745 3166.630 3082.765 ;
        RECT 0.000 3074.715 3165.950 3075.745 ;
        RECT 0.680 3074.635 3165.950 3074.715 ;
        RECT 0.680 3073.565 3166.630 3074.635 ;
        RECT 0.000 3071.495 3166.630 3073.565 ;
        RECT 0.680 3070.345 3166.630 3071.495 ;
        RECT 0.000 3068.275 3166.630 3070.345 ;
        RECT 0.680 3067.125 3166.630 3068.275 ;
        RECT 0.000 3065.735 3166.630 3067.125 ;
        RECT 0.000 3065.515 3165.950 3065.735 ;
        RECT 0.680 3064.625 3165.950 3065.515 ;
        RECT 0.680 3064.365 3166.630 3064.625 ;
        RECT 0.000 3058.265 3166.630 3064.365 ;
        RECT 0.000 3057.115 3165.950 3058.265 ;
        RECT 0.000 3055.505 3166.630 3057.115 ;
        RECT 0.000 3054.355 3165.950 3055.505 ;
        RECT 0.000 3052.285 3166.630 3054.355 ;
        RECT 0.000 3051.135 3165.950 3052.285 ;
        RECT 0.000 3049.610 3166.630 3051.135 ;
        RECT 0.000 3049.065 3166.640 3049.610 ;
        RECT 0.000 3047.915 3165.950 3049.065 ;
        RECT 3166.340 3048.930 3166.640 3049.065 ;
        RECT 3166.030 3048.665 3166.640 3048.930 ;
        RECT 0.000 3042.130 3166.630 3047.915 ;
        RECT 0.000 3039.790 3166.640 3042.130 ;
        RECT 0.000 3038.920 3165.950 3039.790 ;
        RECT 0.680 3038.715 3165.950 3038.920 ;
        RECT 0.680 3037.820 3166.630 3038.715 ;
        RECT 0.000 3037.105 3166.630 3037.820 ;
        RECT 0.000 3035.955 3165.950 3037.105 ;
        RECT 0.000 3033.885 3166.630 3035.955 ;
        RECT 0.000 3032.735 3165.950 3033.885 ;
        RECT 0.000 3030.665 3166.630 3032.735 ;
        RECT 0.000 3029.515 3165.950 3030.665 ;
        RECT 0.000 3028.920 3166.630 3029.515 ;
        RECT 0.680 3027.820 3166.630 3028.920 ;
        RECT 0.000 3018.245 3166.630 3027.820 ;
        RECT 0.000 3017.095 3165.950 3018.245 ;
        RECT 0.000 3015.485 3166.630 3017.095 ;
        RECT 0.000 3014.335 3165.950 3015.485 ;
        RECT 0.000 3012.265 3166.630 3014.335 ;
        RECT 0.000 3011.115 3165.950 3012.265 ;
        RECT 0.000 3009.045 3166.630 3011.115 ;
        RECT 0.000 3007.895 3165.950 3009.045 ;
        RECT 0.000 3006.285 3166.630 3007.895 ;
        RECT 0.000 3005.135 3165.950 3006.285 ;
        RECT 0.000 3003.065 3166.630 3005.135 ;
        RECT 0.000 3001.915 3165.950 3003.065 ;
        RECT 0.000 2997.085 3166.630 3001.915 ;
        RECT 0.000 2995.935 3165.950 2997.085 ;
        RECT 0.000 2993.865 3166.630 2995.935 ;
        RECT 0.000 2992.715 3165.950 2993.865 ;
        RECT 3166.030 2992.870 3166.640 2993.115 ;
        RECT 3166.340 2992.715 3166.640 2992.870 ;
        RECT 0.000 2991.510 3166.640 2992.715 ;
        RECT 0.000 2984.665 3166.630 2991.510 ;
        RECT 0.000 2983.515 3165.950 2984.665 ;
        RECT 0.000 2923.115 3166.630 2983.515 ;
        RECT -0.010 2922.150 0.610 2922.365 ;
        RECT -0.010 2921.965 0.290 2922.150 ;
        RECT 0.680 2921.965 3166.630 2923.115 ;
        RECT -0.010 2921.470 3166.630 2921.965 ;
        RECT 0.000 2913.915 3166.630 2921.470 ;
        RECT 0.680 2912.765 3166.630 2913.915 ;
        RECT 0.000 2910.695 3166.630 2912.765 ;
        RECT 0.680 2909.545 3166.630 2910.695 ;
        RECT 0.000 2904.715 3166.630 2909.545 ;
        RECT -0.010 2903.790 0.610 2903.965 ;
        RECT -0.010 2903.565 0.290 2903.790 ;
        RECT 0.680 2903.565 3166.630 2904.715 ;
        RECT -0.010 2903.110 3166.630 2903.565 ;
        RECT 0.000 2901.495 3166.630 2903.110 ;
        RECT 0.680 2900.345 3166.630 2901.495 ;
        RECT 0.000 2898.735 3166.630 2900.345 ;
        RECT 0.680 2897.585 3166.630 2898.735 ;
        RECT 0.000 2895.515 3166.630 2897.585 ;
        RECT 0.680 2894.365 3166.630 2895.515 ;
        RECT 0.000 2892.295 3166.630 2894.365 ;
        RECT 0.680 2891.145 3166.630 2892.295 ;
        RECT 0.000 2889.535 3166.630 2891.145 ;
        RECT 0.680 2888.385 3166.630 2889.535 ;
        RECT 0.000 2877.115 3166.630 2888.385 ;
        RECT 0.680 2875.965 3166.630 2877.115 ;
        RECT 0.000 2873.895 3166.630 2875.965 ;
        RECT 0.680 2872.745 3166.630 2873.895 ;
        RECT 0.000 2870.675 3166.630 2872.745 ;
        RECT 0.680 2869.525 3166.630 2870.675 ;
        RECT 0.000 2867.915 3166.630 2869.525 ;
        RECT 0.680 2866.765 3166.630 2867.915 ;
        RECT 0.000 2858.715 3166.630 2866.765 ;
        RECT 0.680 2857.565 3166.630 2858.715 ;
        RECT 0.000 2855.495 3166.630 2857.565 ;
        RECT 0.680 2854.345 3166.630 2855.495 ;
        RECT 0.000 2852.275 3166.630 2854.345 ;
        RECT 0.680 2851.125 3166.630 2852.275 ;
        RECT 0.000 2850.745 3166.630 2851.125 ;
        RECT 0.000 2849.635 3165.950 2850.745 ;
        RECT 0.000 2849.515 3166.630 2849.635 ;
        RECT 0.680 2848.365 3166.630 2849.515 ;
        RECT 0.000 2840.735 3166.630 2848.365 ;
        RECT 0.000 2839.625 3165.950 2840.735 ;
        RECT 3166.030 2839.870 3166.640 2840.025 ;
        RECT 3166.340 2839.625 3166.640 2839.870 ;
        RECT 0.000 2839.190 3166.640 2839.625 ;
        RECT 0.000 2833.265 3166.630 2839.190 ;
        RECT 0.000 2832.115 3165.950 2833.265 ;
        RECT 0.000 2830.505 3166.630 2832.115 ;
        RECT 0.000 2829.355 3165.950 2830.505 ;
        RECT 0.000 2827.285 3166.630 2829.355 ;
        RECT 0.000 2826.135 3165.950 2827.285 ;
        RECT 0.000 2825.210 3166.630 2826.135 ;
        RECT 0.000 2824.065 3166.640 2825.210 ;
        RECT 0.000 2823.920 3165.950 2824.065 ;
        RECT 0.680 2822.915 3165.950 2823.920 ;
        RECT 3166.340 2823.850 3166.640 2824.065 ;
        RECT 3166.030 2823.665 3166.640 2823.850 ;
        RECT 0.680 2822.820 3166.630 2822.915 ;
        RECT 0.000 2814.865 3166.630 2822.820 ;
        RECT 0.000 2813.920 3165.950 2814.865 ;
        RECT 0.680 2813.715 3165.950 2813.920 ;
        RECT 0.680 2812.820 3166.630 2813.715 ;
        RECT 0.000 2812.105 3166.630 2812.820 ;
        RECT 0.000 2810.955 3165.950 2812.105 ;
        RECT 0.000 2808.885 3166.630 2810.955 ;
        RECT 0.000 2807.735 3165.950 2808.885 ;
        RECT 0.000 2805.665 3166.630 2807.735 ;
        RECT 0.000 2804.515 3165.950 2805.665 ;
        RECT 0.000 2793.245 3166.630 2804.515 ;
        RECT 0.000 2792.095 3165.950 2793.245 ;
        RECT 0.000 2790.485 3166.630 2792.095 ;
        RECT 0.000 2789.335 3165.950 2790.485 ;
        RECT 0.000 2787.265 3166.630 2789.335 ;
        RECT 0.000 2786.115 3165.950 2787.265 ;
        RECT 0.000 2784.045 3166.630 2786.115 ;
        RECT 0.000 2782.895 3165.950 2784.045 ;
        RECT 0.000 2781.285 3166.630 2782.895 ;
        RECT 0.000 2780.135 3165.950 2781.285 ;
        RECT 0.000 2778.065 3166.630 2780.135 ;
        RECT 0.000 2776.915 3165.950 2778.065 ;
        RECT 0.000 2772.085 3166.630 2776.915 ;
        RECT 0.000 2770.935 3165.950 2772.085 ;
        RECT 0.000 2768.865 3166.630 2770.935 ;
        RECT 0.000 2767.715 3165.950 2768.865 ;
        RECT 0.000 2759.665 3166.630 2767.715 ;
        RECT 0.000 2758.515 3165.950 2759.665 ;
        RECT 0.000 2707.115 3166.630 2758.515 ;
        RECT 0.680 2705.965 3166.630 2707.115 ;
        RECT 0.000 2697.915 3166.630 2705.965 ;
        RECT 0.680 2696.765 3166.630 2697.915 ;
        RECT 0.000 2694.695 3166.630 2696.765 ;
        RECT 0.680 2693.545 3166.630 2694.695 ;
        RECT 0.000 2688.715 3166.630 2693.545 ;
        RECT 0.680 2687.565 3166.630 2688.715 ;
        RECT 0.000 2685.495 3166.630 2687.565 ;
        RECT 0.680 2684.345 3166.630 2685.495 ;
        RECT 0.000 2682.735 3166.630 2684.345 ;
        RECT 0.680 2681.585 3166.630 2682.735 ;
        RECT 0.000 2679.515 3166.630 2681.585 ;
        RECT 0.680 2678.365 3166.630 2679.515 ;
        RECT 0.000 2676.295 3166.630 2678.365 ;
        RECT 0.680 2675.145 3166.630 2676.295 ;
        RECT 0.000 2673.535 3166.630 2675.145 ;
        RECT 0.680 2672.385 3166.630 2673.535 ;
        RECT 0.000 2661.115 3166.630 2672.385 ;
        RECT 0.680 2659.965 3166.630 2661.115 ;
        RECT 0.000 2657.895 3166.630 2659.965 ;
        RECT 0.680 2656.745 3166.630 2657.895 ;
        RECT 0.000 2654.675 3166.630 2656.745 ;
        RECT 0.680 2653.525 3166.630 2654.675 ;
        RECT 0.000 2651.915 3166.630 2653.525 ;
        RECT 0.680 2650.765 3166.630 2651.915 ;
        RECT 0.000 2642.715 3166.630 2650.765 ;
        RECT 0.680 2641.565 3166.630 2642.715 ;
        RECT 0.000 2639.495 3166.630 2641.565 ;
        RECT 0.680 2638.345 3166.630 2639.495 ;
        RECT 0.000 2636.275 3166.630 2638.345 ;
        RECT 0.680 2635.125 3166.630 2636.275 ;
        RECT 0.000 2633.515 3166.630 2635.125 ;
        RECT 0.680 2632.365 3166.630 2633.515 ;
        RECT 0.000 2625.745 3166.630 2632.365 ;
        RECT 0.000 2624.635 3165.950 2625.745 ;
        RECT 0.000 2615.735 3166.630 2624.635 ;
        RECT 0.000 2614.625 3165.950 2615.735 ;
        RECT 0.000 2608.920 3166.630 2614.625 ;
        RECT 0.680 2607.820 3166.630 2608.920 ;
        RECT 0.000 2607.265 3166.630 2607.820 ;
        RECT 0.000 2606.115 3165.950 2607.265 ;
        RECT 0.000 2604.505 3166.630 2606.115 ;
        RECT 0.000 2603.355 3165.950 2604.505 ;
        RECT 0.000 2601.285 3166.630 2603.355 ;
        RECT 0.000 2600.135 3165.950 2601.285 ;
        RECT 0.000 2598.920 3166.630 2600.135 ;
        RECT 0.680 2598.065 3166.630 2598.920 ;
        RECT 0.680 2597.820 3165.950 2598.065 ;
        RECT 0.000 2596.915 3165.950 2597.820 ;
        RECT 0.000 2588.865 3166.630 2596.915 ;
        RECT 0.000 2587.715 3165.950 2588.865 ;
        RECT 0.000 2586.105 3166.630 2587.715 ;
        RECT 0.000 2584.955 3165.950 2586.105 ;
        RECT 0.000 2582.885 3166.630 2584.955 ;
        RECT 0.000 2581.735 3165.950 2582.885 ;
        RECT 0.000 2579.665 3166.630 2581.735 ;
        RECT 0.000 2578.515 3165.950 2579.665 ;
        RECT 3166.030 2578.750 3166.640 2578.915 ;
        RECT 3166.340 2578.515 3166.640 2578.750 ;
        RECT 0.000 2578.070 3166.640 2578.515 ;
        RECT 0.000 2567.245 3166.630 2578.070 ;
        RECT 0.000 2566.095 3165.950 2567.245 ;
        RECT 0.000 2564.485 3166.630 2566.095 ;
        RECT 0.000 2563.335 3165.950 2564.485 ;
        RECT 0.000 2561.265 3166.630 2563.335 ;
        RECT 0.000 2560.115 3165.950 2561.265 ;
        RECT 0.000 2558.045 3166.630 2560.115 ;
        RECT 0.000 2556.895 3165.950 2558.045 ;
        RECT 0.000 2555.285 3166.630 2556.895 ;
        RECT 0.000 2554.135 3165.950 2555.285 ;
        RECT 0.000 2552.065 3166.630 2554.135 ;
        RECT 0.000 2550.915 3165.950 2552.065 ;
        RECT 0.000 2546.085 3166.630 2550.915 ;
        RECT 0.000 2544.935 3165.950 2546.085 ;
        RECT 0.000 2542.865 3166.630 2544.935 ;
        RECT 0.000 2541.715 3165.950 2542.865 ;
        RECT 0.000 2533.665 3166.630 2541.715 ;
        RECT 0.000 2532.515 3165.950 2533.665 ;
        RECT 0.000 2491.115 3166.630 2532.515 ;
        RECT 0.680 2489.965 3166.630 2491.115 ;
        RECT 0.000 2481.915 3166.630 2489.965 ;
        RECT 0.680 2480.765 3166.630 2481.915 ;
        RECT 0.000 2478.695 3166.630 2480.765 ;
        RECT 0.680 2477.545 3166.630 2478.695 ;
        RECT 0.000 2472.715 3166.630 2477.545 ;
        RECT 0.680 2471.565 3166.630 2472.715 ;
        RECT 0.000 2469.495 3166.630 2471.565 ;
        RECT 0.680 2468.345 3166.630 2469.495 ;
        RECT 0.000 2466.735 3166.630 2468.345 ;
        RECT 0.680 2465.585 3166.630 2466.735 ;
        RECT 0.000 2463.515 3166.630 2465.585 ;
        RECT 0.680 2462.365 3166.630 2463.515 ;
        RECT 0.000 2460.295 3166.630 2462.365 ;
        RECT 0.680 2459.145 3166.630 2460.295 ;
        RECT 0.000 2458.010 3166.630 2459.145 ;
        RECT -0.010 2457.535 3166.630 2458.010 ;
        RECT -0.010 2457.330 0.290 2457.535 ;
        RECT -0.010 2457.135 0.610 2457.330 ;
        RECT 0.680 2456.385 3166.630 2457.535 ;
        RECT 0.000 2445.115 3166.630 2456.385 ;
        RECT 0.680 2443.965 3166.630 2445.115 ;
        RECT 0.000 2442.370 3166.630 2443.965 ;
        RECT -0.010 2441.895 3166.630 2442.370 ;
        RECT -0.010 2441.690 0.290 2441.895 ;
        RECT -0.010 2441.495 0.610 2441.690 ;
        RECT 0.680 2440.745 3166.630 2441.895 ;
        RECT 0.000 2438.675 3166.630 2440.745 ;
        RECT 0.680 2437.525 3166.630 2438.675 ;
        RECT 0.000 2435.915 3166.630 2437.525 ;
        RECT 0.680 2434.765 3166.630 2435.915 ;
        RECT 0.000 2426.715 3166.630 2434.765 ;
        RECT 0.680 2425.565 3166.630 2426.715 ;
        RECT 0.000 2423.495 3166.630 2425.565 ;
        RECT 0.680 2422.345 3166.630 2423.495 ;
        RECT 0.000 2420.275 3166.630 2422.345 ;
        RECT 0.680 2419.125 3166.630 2420.275 ;
        RECT 0.000 2417.515 3166.630 2419.125 ;
        RECT 0.680 2416.365 3166.630 2417.515 ;
        RECT 0.000 2393.920 3166.630 2416.365 ;
        RECT 0.680 2392.820 3166.630 2393.920 ;
        RECT 0.000 2383.920 3166.630 2392.820 ;
        RECT 0.680 2382.820 3166.630 2383.920 ;
        RECT 0.000 2162.815 3166.630 2382.820 ;
        RECT 0.000 2088.615 3122.620 2162.815 ;
      LAYER met3 ;
        RECT 3122.620 2088.615 3167.855 2162.815 ;
      LAYER met3 ;
        RECT 0.000 1853.115 3166.630 2088.615 ;
        RECT 0.680 1851.965 3166.630 1853.115 ;
        RECT 0.000 1843.915 3166.630 1851.965 ;
        RECT -0.010 1842.990 0.610 1843.165 ;
        RECT -0.010 1842.765 0.290 1842.990 ;
        RECT 0.680 1842.765 3166.630 1843.915 ;
        RECT -0.010 1842.310 3166.630 1842.765 ;
        RECT 0.000 1840.695 3166.630 1842.310 ;
        RECT 0.680 1839.545 3166.630 1840.695 ;
        RECT 0.000 1834.715 3166.630 1839.545 ;
        RECT 0.680 1833.565 3166.630 1834.715 ;
        RECT 0.000 1831.495 3166.630 1833.565 ;
        RECT 0.680 1830.345 3166.630 1831.495 ;
        RECT 0.000 1828.735 3166.630 1830.345 ;
        RECT 0.680 1827.585 3166.630 1828.735 ;
        RECT 0.000 1825.515 3166.630 1827.585 ;
        RECT 0.680 1824.365 3166.630 1825.515 ;
        RECT 0.000 1822.295 3166.630 1824.365 ;
        RECT 0.680 1821.145 3166.630 1822.295 ;
        RECT 0.000 1819.535 3166.630 1821.145 ;
        RECT 0.680 1818.385 3166.630 1819.535 ;
        RECT 0.000 1807.115 3166.630 1818.385 ;
        RECT 0.680 1805.965 3166.630 1807.115 ;
        RECT 0.000 1803.895 3166.630 1805.965 ;
        RECT 0.680 1802.745 3166.630 1803.895 ;
        RECT 0.000 1800.675 3166.630 1802.745 ;
        RECT 0.680 1799.525 3166.630 1800.675 ;
        RECT 0.000 1797.915 3166.630 1799.525 ;
        RECT 0.680 1796.765 3166.630 1797.915 ;
        RECT 0.000 1788.715 3166.630 1796.765 ;
        RECT 0.680 1787.565 3166.630 1788.715 ;
        RECT 0.000 1785.495 3166.630 1787.565 ;
        RECT 0.680 1784.345 3166.630 1785.495 ;
        RECT 0.000 1782.275 3166.630 1784.345 ;
        RECT 0.680 1781.125 3166.630 1782.275 ;
        RECT 0.000 1779.515 3166.630 1781.125 ;
        RECT 0.680 1778.365 3166.630 1779.515 ;
        RECT 0.000 1749.450 3166.630 1778.365 ;
        RECT -0.010 1748.920 3166.630 1749.450 ;
        RECT -0.010 1748.770 0.290 1748.920 ;
        RECT -0.010 1748.520 0.610 1748.770 ;
        RECT 0.680 1747.820 3166.630 1748.920 ;
        RECT 0.000 1741.290 3166.630 1747.820 ;
        RECT 0.000 1740.745 3166.640 1741.290 ;
        RECT 0.000 1739.635 3165.950 1740.745 ;
        RECT 3166.340 1740.610 3166.640 1740.745 ;
        RECT 3166.030 1740.345 3166.640 1740.610 ;
        RECT 0.000 1738.920 3166.630 1739.635 ;
        RECT 0.680 1737.820 3166.630 1738.920 ;
        RECT 0.000 1730.735 3166.630 1737.820 ;
        RECT 0.000 1729.625 3165.950 1730.735 ;
        RECT 0.000 1721.265 3166.630 1729.625 ;
        RECT 0.000 1720.115 3165.950 1721.265 ;
        RECT 0.000 1718.505 3166.630 1720.115 ;
        RECT 0.000 1717.355 3165.950 1718.505 ;
        RECT 0.000 1715.285 3166.630 1717.355 ;
        RECT 0.000 1714.135 3165.950 1715.285 ;
        RECT 0.000 1712.065 3166.630 1714.135 ;
        RECT 0.000 1710.915 3165.950 1712.065 ;
        RECT 0.000 1702.865 3166.630 1710.915 ;
        RECT 0.000 1701.715 3165.950 1702.865 ;
        RECT 0.000 1700.105 3166.630 1701.715 ;
        RECT 0.000 1698.955 3165.950 1700.105 ;
        RECT 0.000 1696.885 3166.630 1698.955 ;
        RECT 0.000 1695.735 3165.950 1696.885 ;
        RECT 0.000 1693.665 3166.630 1695.735 ;
        RECT 0.000 1692.515 3165.950 1693.665 ;
        RECT 3166.030 1692.710 3166.640 1692.915 ;
        RECT 3166.340 1692.515 3166.640 1692.710 ;
        RECT 0.000 1690.670 3166.640 1692.515 ;
        RECT 0.000 1681.245 3166.630 1690.670 ;
        RECT 0.000 1680.095 3165.950 1681.245 ;
        RECT 0.000 1678.485 3166.630 1680.095 ;
        RECT 0.000 1677.335 3165.950 1678.485 ;
        RECT 0.000 1675.265 3166.630 1677.335 ;
        RECT 0.000 1674.115 3165.950 1675.265 ;
        RECT 3166.030 1674.350 3166.640 1674.515 ;
        RECT 3166.340 1674.115 3166.640 1674.350 ;
        RECT 0.000 1672.990 3166.640 1674.115 ;
        RECT 0.000 1672.045 3166.630 1672.990 ;
        RECT 0.000 1670.895 3165.950 1672.045 ;
        RECT 0.000 1669.285 3166.630 1670.895 ;
        RECT 0.000 1668.135 3165.950 1669.285 ;
        RECT 0.000 1666.065 3166.630 1668.135 ;
        RECT 0.000 1664.915 3165.950 1666.065 ;
        RECT 0.000 1660.085 3166.630 1664.915 ;
        RECT 0.000 1658.935 3165.950 1660.085 ;
        RECT 0.000 1656.865 3166.630 1658.935 ;
        RECT 0.000 1655.715 3165.950 1656.865 ;
        RECT 0.000 1648.810 3166.630 1655.715 ;
        RECT 0.000 1647.665 3166.640 1648.810 ;
        RECT 0.000 1646.515 3165.950 1647.665 ;
        RECT 3166.340 1647.450 3166.640 1647.665 ;
        RECT 3166.030 1647.265 3166.640 1647.450 ;
        RECT 0.000 1637.115 3166.630 1646.515 ;
        RECT 0.680 1635.965 3166.630 1637.115 ;
        RECT 0.000 1627.915 3166.630 1635.965 ;
        RECT 0.680 1626.765 3166.630 1627.915 ;
        RECT 0.000 1624.695 3166.630 1626.765 ;
        RECT 0.680 1623.545 3166.630 1624.695 ;
        RECT 0.000 1618.715 3166.630 1623.545 ;
        RECT 0.680 1617.565 3166.630 1618.715 ;
        RECT 0.000 1615.495 3166.630 1617.565 ;
        RECT 0.680 1614.345 3166.630 1615.495 ;
        RECT 0.000 1612.735 3166.630 1614.345 ;
        RECT 0.680 1611.585 3166.630 1612.735 ;
        RECT 0.000 1610.050 3166.630 1611.585 ;
        RECT -0.010 1609.515 3166.630 1610.050 ;
        RECT -0.010 1609.370 0.290 1609.515 ;
        RECT -0.010 1609.115 0.610 1609.370 ;
        RECT 0.680 1608.365 3166.630 1609.515 ;
        RECT 0.000 1606.295 3166.630 1608.365 ;
        RECT 0.680 1605.145 3166.630 1606.295 ;
        RECT 0.000 1603.535 3166.630 1605.145 ;
        RECT 0.680 1602.385 3166.630 1603.535 ;
        RECT 0.000 1591.115 3166.630 1602.385 ;
        RECT 0.680 1589.965 3166.630 1591.115 ;
        RECT 0.000 1587.895 3166.630 1589.965 ;
        RECT 0.680 1586.745 3166.630 1587.895 ;
        RECT 0.000 1584.675 3166.630 1586.745 ;
        RECT 0.680 1583.525 3166.630 1584.675 ;
        RECT 0.000 1581.915 3166.630 1583.525 ;
        RECT 0.680 1580.765 3166.630 1581.915 ;
        RECT 0.000 1572.715 3166.630 1580.765 ;
        RECT 0.680 1571.565 3166.630 1572.715 ;
        RECT 0.000 1569.495 3166.630 1571.565 ;
        RECT 0.680 1568.345 3166.630 1569.495 ;
        RECT 0.000 1566.275 3166.630 1568.345 ;
        RECT 0.680 1565.125 3166.630 1566.275 ;
        RECT 0.000 1563.515 3166.630 1565.125 ;
        RECT 0.680 1562.365 3166.630 1563.515 ;
        RECT 0.000 1533.920 3166.630 1562.365 ;
        RECT 0.680 1532.820 3166.630 1533.920 ;
        RECT 0.000 1524.370 3166.630 1532.820 ;
        RECT -0.010 1523.920 3166.630 1524.370 ;
        RECT -0.010 1523.690 0.290 1523.920 ;
        RECT -0.010 1523.520 0.610 1523.690 ;
        RECT 0.680 1522.820 3166.630 1523.920 ;
        RECT 0.000 1515.745 3166.630 1522.820 ;
        RECT 0.000 1514.635 3165.950 1515.745 ;
        RECT 0.000 1505.735 3166.630 1514.635 ;
        RECT 0.000 1504.625 3165.950 1505.735 ;
        RECT 0.000 1495.265 3166.630 1504.625 ;
        RECT 0.000 1494.115 3165.950 1495.265 ;
        RECT 0.000 1492.505 3166.630 1494.115 ;
        RECT 0.000 1491.355 3165.950 1492.505 ;
        RECT 0.000 1489.285 3166.630 1491.355 ;
        RECT 0.000 1488.135 3165.950 1489.285 ;
        RECT 0.000 1486.065 3166.630 1488.135 ;
        RECT 0.000 1484.915 3165.950 1486.065 ;
        RECT 0.000 1476.865 3166.630 1484.915 ;
        RECT 0.000 1475.715 3165.950 1476.865 ;
        RECT 0.000 1474.105 3166.630 1475.715 ;
        RECT 0.000 1472.955 3165.950 1474.105 ;
        RECT 0.000 1471.330 3166.630 1472.955 ;
        RECT 0.000 1470.885 3166.640 1471.330 ;
        RECT 0.000 1469.735 3165.950 1470.885 ;
        RECT 3166.340 1470.650 3166.640 1470.885 ;
        RECT 3166.030 1470.485 3166.640 1470.650 ;
        RECT 0.000 1467.665 3166.630 1469.735 ;
        RECT 0.000 1466.515 3165.950 1467.665 ;
        RECT 0.000 1455.690 3166.630 1466.515 ;
        RECT 0.000 1455.245 3166.640 1455.690 ;
        RECT 0.000 1454.095 3165.950 1455.245 ;
        RECT 3166.340 1455.010 3166.640 1455.245 ;
        RECT 3166.030 1454.845 3166.640 1455.010 ;
        RECT 0.000 1452.485 3166.630 1454.095 ;
        RECT 0.000 1451.335 3165.950 1452.485 ;
        RECT 0.000 1449.265 3166.630 1451.335 ;
        RECT 0.000 1448.115 3165.950 1449.265 ;
        RECT 0.000 1446.045 3166.630 1448.115 ;
        RECT 0.000 1444.895 3165.950 1446.045 ;
        RECT 0.000 1443.285 3166.630 1444.895 ;
        RECT 0.000 1442.135 3165.950 1443.285 ;
        RECT 0.000 1440.065 3166.630 1442.135 ;
        RECT 0.000 1438.915 3165.950 1440.065 ;
        RECT 3166.030 1439.070 3166.640 1439.315 ;
        RECT 3166.340 1438.915 3166.640 1439.070 ;
        RECT 0.000 1438.390 3166.640 1438.915 ;
        RECT 0.000 1434.085 3166.630 1438.390 ;
        RECT 0.000 1432.935 3165.950 1434.085 ;
        RECT 0.000 1430.865 3166.630 1432.935 ;
        RECT 0.000 1429.715 3165.950 1430.865 ;
        RECT 0.000 1421.665 3166.630 1429.715 ;
        RECT 0.000 1421.115 3165.950 1421.665 ;
        RECT 0.680 1420.515 3165.950 1421.115 ;
        RECT 0.680 1419.965 3166.630 1420.515 ;
        RECT 0.000 1411.915 3166.630 1419.965 ;
        RECT 0.680 1410.765 3166.630 1411.915 ;
        RECT 0.000 1408.695 3166.630 1410.765 ;
        RECT 0.680 1407.545 3166.630 1408.695 ;
        RECT 0.000 1402.715 3166.630 1407.545 ;
        RECT 0.680 1401.565 3166.630 1402.715 ;
        RECT 0.000 1399.495 3166.630 1401.565 ;
        RECT 0.680 1398.345 3166.630 1399.495 ;
        RECT 0.000 1397.210 3166.630 1398.345 ;
        RECT -0.010 1396.735 3166.630 1397.210 ;
        RECT -0.010 1396.530 0.290 1396.735 ;
        RECT -0.010 1396.335 0.610 1396.530 ;
        RECT 0.680 1395.585 3166.630 1396.735 ;
        RECT 0.000 1393.515 3166.630 1395.585 ;
        RECT 0.680 1392.365 3166.630 1393.515 ;
        RECT 0.000 1390.295 3166.630 1392.365 ;
        RECT 0.680 1389.145 3166.630 1390.295 ;
        RECT 0.000 1387.535 3166.630 1389.145 ;
        RECT 0.680 1386.385 3166.630 1387.535 ;
        RECT 0.000 1375.115 3166.630 1386.385 ;
        RECT 0.680 1373.965 3166.630 1375.115 ;
        RECT 0.000 1371.895 3166.630 1373.965 ;
        RECT 0.680 1370.745 3166.630 1371.895 ;
        RECT 0.000 1368.675 3166.630 1370.745 ;
        RECT 0.680 1367.525 3166.630 1368.675 ;
        RECT 0.000 1365.915 3166.630 1367.525 ;
        RECT 0.680 1364.765 3166.630 1365.915 ;
        RECT 0.000 1356.715 3166.630 1364.765 ;
        RECT 0.680 1355.565 3166.630 1356.715 ;
        RECT 0.000 1353.495 3166.630 1355.565 ;
        RECT 0.680 1352.345 3166.630 1353.495 ;
        RECT 0.000 1350.275 3166.630 1352.345 ;
        RECT 0.680 1349.125 3166.630 1350.275 ;
        RECT 0.000 1347.515 3166.630 1349.125 ;
        RECT 0.680 1346.365 3166.630 1347.515 ;
        RECT 0.000 1318.920 3166.630 1346.365 ;
        RECT 0.680 1317.820 3166.630 1318.920 ;
        RECT 0.000 1308.920 3166.630 1317.820 ;
        RECT 0.680 1307.820 3166.630 1308.920 ;
        RECT 0.000 1290.745 3166.630 1307.820 ;
        RECT 0.000 1289.635 3165.950 1290.745 ;
        RECT 0.000 1280.735 3166.630 1289.635 ;
        RECT 0.000 1279.625 3165.950 1280.735 ;
        RECT 0.000 1270.265 3166.630 1279.625 ;
        RECT 0.000 1269.115 3165.950 1270.265 ;
        RECT 0.000 1268.010 3166.630 1269.115 ;
        RECT 0.000 1267.505 3166.640 1268.010 ;
        RECT 0.000 1266.355 3165.950 1267.505 ;
        RECT 3166.340 1267.330 3166.640 1267.505 ;
        RECT 3166.030 1267.105 3166.640 1267.330 ;
        RECT 0.000 1264.285 3166.630 1266.355 ;
        RECT 0.000 1263.135 3165.950 1264.285 ;
        RECT 0.000 1261.065 3166.630 1263.135 ;
        RECT 0.000 1259.915 3165.950 1261.065 ;
        RECT 0.000 1251.865 3166.630 1259.915 ;
        RECT 0.000 1250.715 3165.950 1251.865 ;
        RECT 0.000 1249.105 3166.630 1250.715 ;
        RECT 0.000 1247.955 3165.950 1249.105 ;
        RECT 0.000 1245.885 3166.630 1247.955 ;
        RECT 0.000 1244.735 3165.950 1245.885 ;
        RECT 0.000 1242.665 3166.630 1244.735 ;
        RECT 0.000 1241.515 3165.950 1242.665 ;
        RECT 0.000 1230.245 3166.630 1241.515 ;
        RECT 0.000 1229.095 3165.950 1230.245 ;
        RECT 0.000 1227.485 3166.630 1229.095 ;
        RECT 0.000 1226.335 3165.950 1227.485 ;
        RECT 0.000 1224.265 3166.630 1226.335 ;
        RECT 0.000 1223.115 3165.950 1224.265 ;
        RECT 0.000 1221.045 3166.630 1223.115 ;
        RECT 0.000 1219.895 3165.950 1221.045 ;
        RECT 0.000 1218.285 3166.630 1219.895 ;
        RECT 0.000 1217.135 3165.950 1218.285 ;
        RECT 0.000 1215.065 3166.630 1217.135 ;
        RECT 0.000 1213.915 3165.950 1215.065 ;
        RECT 0.000 1209.085 3166.630 1213.915 ;
        RECT 0.000 1207.935 3165.950 1209.085 ;
        RECT 0.000 1205.865 3166.630 1207.935 ;
        RECT 0.000 1205.115 3165.950 1205.865 ;
        RECT 0.680 1204.715 3165.950 1205.115 ;
        RECT 0.680 1203.965 3166.630 1204.715 ;
        RECT 0.000 1196.665 3166.630 1203.965 ;
        RECT 0.000 1195.915 3165.950 1196.665 ;
        RECT 0.680 1195.515 3165.950 1195.915 ;
        RECT 0.680 1194.765 3166.630 1195.515 ;
        RECT 0.000 1192.695 3166.630 1194.765 ;
        RECT 0.680 1191.545 3166.630 1192.695 ;
        RECT 0.000 1186.715 3166.630 1191.545 ;
        RECT 0.680 1185.565 3166.630 1186.715 ;
        RECT 0.000 1183.495 3166.630 1185.565 ;
        RECT 0.680 1182.345 3166.630 1183.495 ;
        RECT 0.000 1180.735 3166.630 1182.345 ;
        RECT 0.680 1179.585 3166.630 1180.735 ;
        RECT 0.000 1177.515 3166.630 1179.585 ;
        RECT -0.010 1176.590 0.610 1176.765 ;
        RECT -0.010 1176.365 0.290 1176.590 ;
        RECT 0.680 1176.365 3166.630 1177.515 ;
        RECT -0.010 1175.910 3166.630 1176.365 ;
        RECT 0.000 1174.850 3166.630 1175.910 ;
        RECT -0.010 1174.295 3166.630 1174.850 ;
        RECT -0.010 1174.170 0.290 1174.295 ;
        RECT -0.010 1173.895 0.610 1174.170 ;
        RECT 0.680 1173.145 3166.630 1174.295 ;
        RECT 0.000 1171.535 3166.630 1173.145 ;
        RECT 0.680 1170.385 3166.630 1171.535 ;
        RECT 0.000 1159.115 3166.630 1170.385 ;
        RECT 0.680 1157.965 3166.630 1159.115 ;
        RECT 0.000 1155.895 3166.630 1157.965 ;
        RECT 0.680 1154.745 3166.630 1155.895 ;
        RECT 0.000 1152.675 3166.630 1154.745 ;
        RECT 0.680 1151.525 3166.630 1152.675 ;
        RECT 0.000 1150.370 3166.630 1151.525 ;
        RECT -0.010 1149.915 3166.630 1150.370 ;
        RECT -0.010 1149.690 0.290 1149.915 ;
        RECT -0.010 1149.515 0.610 1149.690 ;
        RECT 0.680 1148.765 3166.630 1149.915 ;
        RECT 0.000 1140.715 3166.630 1148.765 ;
        RECT 0.680 1139.565 3166.630 1140.715 ;
        RECT 0.000 1137.495 3166.630 1139.565 ;
        RECT 0.680 1136.345 3166.630 1137.495 ;
        RECT 0.000 1134.275 3166.630 1136.345 ;
        RECT 0.680 1133.125 3166.630 1134.275 ;
        RECT 0.000 1131.515 3166.630 1133.125 ;
        RECT 0.680 1130.365 3166.630 1131.515 ;
        RECT 0.000 1103.920 3166.630 1130.365 ;
        RECT 0.680 1102.820 3166.630 1103.920 ;
        RECT 0.000 1093.920 3166.630 1102.820 ;
        RECT 0.680 1092.820 3166.630 1093.920 ;
        RECT 0.000 1065.745 3166.630 1092.820 ;
        RECT 0.000 1064.635 3165.950 1065.745 ;
        RECT 0.000 1055.735 3166.630 1064.635 ;
        RECT 0.000 1054.625 3165.950 1055.735 ;
        RECT 0.000 1045.265 3166.630 1054.625 ;
        RECT 0.000 1044.115 3165.950 1045.265 ;
        RECT 0.000 1042.505 3166.630 1044.115 ;
        RECT 0.000 1041.355 3165.950 1042.505 ;
        RECT 0.000 1039.285 3166.630 1041.355 ;
        RECT 0.000 1038.135 3165.950 1039.285 ;
        RECT 0.000 1036.065 3166.630 1038.135 ;
        RECT 0.000 1034.915 3165.950 1036.065 ;
        RECT 0.000 1026.865 3166.630 1034.915 ;
        RECT 0.000 1025.715 3165.950 1026.865 ;
        RECT 0.000 1024.570 3166.630 1025.715 ;
        RECT 0.000 1024.105 3166.640 1024.570 ;
        RECT 0.000 1022.955 3165.950 1024.105 ;
        RECT 3166.340 1023.890 3166.640 1024.105 ;
        RECT 3166.030 1023.705 3166.640 1023.890 ;
        RECT 0.000 1020.885 3166.630 1022.955 ;
        RECT 0.000 1019.735 3165.950 1020.885 ;
        RECT 0.000 1017.665 3166.630 1019.735 ;
        RECT 0.000 1016.515 3165.950 1017.665 ;
        RECT 0.000 1005.245 3166.630 1016.515 ;
        RECT 0.000 1004.095 3165.950 1005.245 ;
        RECT 0.000 1002.485 3166.630 1004.095 ;
        RECT 0.000 1001.335 3165.950 1002.485 ;
        RECT 0.000 999.265 3166.630 1001.335 ;
        RECT 0.000 998.115 3165.950 999.265 ;
        RECT 0.000 996.045 3166.630 998.115 ;
        RECT 0.000 994.895 3165.950 996.045 ;
        RECT 3166.030 995.030 3166.640 995.295 ;
        RECT 3166.340 994.895 3166.640 995.030 ;
        RECT 0.000 993.670 3166.640 994.895 ;
        RECT 0.000 993.285 3166.630 993.670 ;
        RECT 0.000 992.135 3165.950 993.285 ;
        RECT 0.000 990.065 3166.630 992.135 ;
        RECT 0.000 989.120 3165.950 990.065 ;
        RECT 0.680 988.915 3165.950 989.120 ;
        RECT 0.680 987.960 3166.630 988.915 ;
        RECT 0.000 984.085 3166.630 987.960 ;
        RECT 0.000 982.935 3165.950 984.085 ;
        RECT 0.000 980.865 3166.630 982.935 ;
        RECT 0.000 979.920 3165.950 980.865 ;
        RECT 0.680 979.715 3165.950 979.920 ;
        RECT 0.680 978.760 3166.630 979.715 ;
        RECT 0.000 976.700 3166.630 978.760 ;
        RECT 0.680 975.540 3166.630 976.700 ;
        RECT 0.000 971.665 3166.630 975.540 ;
        RECT 0.000 970.720 3165.950 971.665 ;
        RECT 0.680 970.515 3165.950 970.720 ;
        RECT 0.680 969.560 3166.630 970.515 ;
        RECT 0.000 967.500 3166.630 969.560 ;
        RECT 0.680 966.340 3166.630 967.500 ;
        RECT 0.000 964.740 3166.630 966.340 ;
        RECT 0.680 963.580 3166.630 964.740 ;
        RECT 0.000 962.010 3166.630 963.580 ;
        RECT -0.010 961.520 3166.630 962.010 ;
        RECT -0.010 961.330 0.290 961.520 ;
        RECT -0.010 961.120 0.610 961.330 ;
        RECT 0.680 960.360 3166.630 961.520 ;
        RECT 0.000 958.300 3166.630 960.360 ;
        RECT 0.680 957.140 3166.630 958.300 ;
        RECT 0.000 955.540 3166.630 957.140 ;
        RECT 0.680 954.380 3166.630 955.540 ;
        RECT 0.000 944.330 3166.630 954.380 ;
        RECT -0.010 943.120 3166.630 944.330 ;
        RECT -0.010 942.970 0.290 943.120 ;
        RECT -0.010 942.720 0.610 942.970 ;
        RECT 0.680 941.960 3166.630 943.120 ;
        RECT 0.000 939.900 3166.630 941.960 ;
        RECT 0.680 938.740 3166.630 939.900 ;
        RECT 0.000 936.680 3166.630 938.740 ;
        RECT 0.680 935.520 3166.630 936.680 ;
        RECT 0.000 933.920 3166.630 935.520 ;
        RECT 0.680 932.760 3166.630 933.920 ;
        RECT 0.000 924.720 3166.630 932.760 ;
        RECT 0.680 923.560 3166.630 924.720 ;
        RECT 0.000 921.500 3166.630 923.560 ;
        RECT 0.680 920.340 3166.630 921.500 ;
        RECT 0.000 918.280 3166.630 920.340 ;
        RECT 0.680 917.120 3166.630 918.280 ;
        RECT 0.000 915.520 3166.630 917.120 ;
        RECT 0.680 914.360 3166.630 915.520 ;
        RECT 0.000 889.930 3166.630 914.360 ;
        RECT -0.010 888.950 3166.630 889.930 ;
        RECT 0.000 888.920 3166.630 888.950 ;
        RECT 0.680 887.820 3166.630 888.920 ;
        RECT 0.000 878.920 3166.630 887.820 ;
        RECT 0.680 877.820 3166.630 878.920 ;
        RECT 0.000 840.745 3166.630 877.820 ;
        RECT 0.000 839.635 3165.950 840.745 ;
        RECT 0.000 830.735 3166.630 839.635 ;
        RECT 0.000 829.625 3165.950 830.735 ;
        RECT 0.000 819.265 3166.630 829.625 ;
        RECT 0.000 818.115 3165.950 819.265 ;
        RECT 0.000 816.505 3166.630 818.115 ;
        RECT 0.000 815.355 3165.950 816.505 ;
        RECT 0.000 813.285 3166.630 815.355 ;
        RECT 0.000 812.135 3165.950 813.285 ;
        RECT 0.000 810.065 3166.630 812.135 ;
        RECT 0.000 808.915 3165.950 810.065 ;
        RECT 0.000 800.865 3166.630 808.915 ;
        RECT 0.000 799.715 3165.950 800.865 ;
        RECT 0.000 798.105 3166.630 799.715 ;
        RECT 0.000 796.955 3165.950 798.105 ;
        RECT 3166.030 797.150 3166.640 797.355 ;
        RECT 3166.340 796.955 3166.640 797.150 ;
        RECT 0.000 796.470 3166.640 796.955 ;
        RECT 0.000 794.885 3166.630 796.470 ;
        RECT 0.000 793.735 3165.950 794.885 ;
        RECT 0.000 791.665 3166.630 793.735 ;
        RECT 0.000 790.515 3165.950 791.665 ;
        RECT 0.000 779.245 3166.630 790.515 ;
        RECT 0.000 778.095 3165.950 779.245 ;
        RECT 0.000 776.485 3166.630 778.095 ;
        RECT 0.000 775.335 3165.950 776.485 ;
        RECT 0.000 773.265 3166.630 775.335 ;
        RECT 0.000 773.120 3165.950 773.265 ;
        RECT 0.680 772.115 3165.950 773.120 ;
        RECT 0.680 771.960 3166.630 772.115 ;
        RECT 0.000 770.045 3166.630 771.960 ;
        RECT 0.000 768.895 3165.950 770.045 ;
        RECT 0.000 767.285 3166.630 768.895 ;
        RECT 0.000 766.135 3165.950 767.285 ;
        RECT 0.000 764.065 3166.630 766.135 ;
        RECT 0.000 763.920 3165.950 764.065 ;
        RECT 0.680 762.915 3165.950 763.920 ;
        RECT 0.680 762.760 3166.630 762.915 ;
        RECT 0.000 760.700 3166.630 762.760 ;
        RECT 0.680 759.540 3166.630 760.700 ;
        RECT 0.000 758.085 3166.630 759.540 ;
        RECT 0.000 756.935 3165.950 758.085 ;
        RECT 0.000 754.865 3166.630 756.935 ;
        RECT 0.000 754.720 3165.950 754.865 ;
        RECT 0.680 753.715 3165.950 754.720 ;
        RECT 0.680 753.560 3166.630 753.715 ;
        RECT 0.000 751.500 3166.630 753.560 ;
        RECT 0.680 750.340 3166.630 751.500 ;
        RECT 0.000 748.740 3166.630 750.340 ;
        RECT 0.680 747.580 3166.630 748.740 ;
        RECT 0.000 745.665 3166.630 747.580 ;
        RECT 0.000 745.520 3165.950 745.665 ;
        RECT 0.680 744.515 3165.950 745.520 ;
        RECT 0.680 744.360 3166.630 744.515 ;
        RECT 0.000 742.300 3166.630 744.360 ;
        RECT 0.680 741.140 3166.630 742.300 ;
        RECT 0.000 739.540 3166.630 741.140 ;
        RECT 0.680 738.380 3166.630 739.540 ;
        RECT 0.000 727.120 3166.630 738.380 ;
        RECT 0.680 725.960 3166.630 727.120 ;
        RECT 0.000 723.900 3166.630 725.960 ;
        RECT 0.680 722.740 3166.630 723.900 ;
        RECT 0.000 720.680 3166.630 722.740 ;
        RECT 0.680 719.520 3166.630 720.680 ;
        RECT 0.000 717.920 3166.630 719.520 ;
        RECT 0.680 716.760 3166.630 717.920 ;
        RECT 0.000 708.720 3166.630 716.760 ;
        RECT 0.680 707.560 3166.630 708.720 ;
        RECT 0.000 705.500 3166.630 707.560 ;
        RECT 0.680 704.340 3166.630 705.500 ;
        RECT 0.000 702.280 3166.630 704.340 ;
        RECT 0.680 701.120 3166.630 702.280 ;
        RECT 0.000 699.520 3166.630 701.120 ;
        RECT 0.680 698.360 3166.630 699.520 ;
        RECT 0.000 675.050 3166.630 698.360 ;
        RECT -0.010 673.920 3166.630 675.050 ;
        RECT -0.010 673.690 0.290 673.920 ;
        RECT -0.010 673.520 0.610 673.690 ;
        RECT 0.680 672.820 3166.630 673.920 ;
        RECT 0.000 663.920 3166.630 672.820 ;
        RECT 0.680 662.820 3166.630 663.920 ;
        RECT 0.000 615.745 3166.630 662.820 ;
        RECT 0.000 614.635 3165.950 615.745 ;
        RECT 0.000 605.735 3166.630 614.635 ;
        RECT 0.000 604.625 3165.950 605.735 ;
        RECT 0.000 594.265 3166.630 604.625 ;
        RECT 0.000 593.115 3165.950 594.265 ;
        RECT 0.000 591.505 3166.630 593.115 ;
        RECT 0.000 590.355 3165.950 591.505 ;
        RECT 0.000 588.285 3166.630 590.355 ;
        RECT 0.000 587.135 3165.950 588.285 ;
        RECT 0.000 585.065 3166.630 587.135 ;
        RECT 0.000 583.915 3165.950 585.065 ;
        RECT 0.000 575.865 3166.630 583.915 ;
        RECT 0.000 574.715 3165.950 575.865 ;
        RECT 0.000 573.105 3166.630 574.715 ;
        RECT 0.000 571.955 3165.950 573.105 ;
        RECT 0.000 569.885 3166.630 571.955 ;
        RECT 0.000 568.735 3165.950 569.885 ;
        RECT 0.000 566.665 3166.630 568.735 ;
        RECT 0.000 565.515 3165.950 566.665 ;
        RECT 0.000 554.690 3166.630 565.515 ;
        RECT 0.000 554.245 3166.640 554.690 ;
        RECT 0.000 553.095 3165.950 554.245 ;
        RECT 3166.340 554.010 3166.640 554.245 ;
        RECT 3166.030 553.845 3166.640 554.010 ;
        RECT 0.000 551.485 3166.630 553.095 ;
        RECT 0.000 550.335 3165.950 551.485 ;
        RECT 0.000 548.265 3166.630 550.335 ;
        RECT 0.000 547.115 3165.950 548.265 ;
        RECT 0.000 545.045 3166.630 547.115 ;
        RECT 0.000 543.895 3165.950 545.045 ;
        RECT 0.000 542.285 3166.630 543.895 ;
        RECT 0.000 541.135 3165.950 542.285 ;
        RECT 0.000 539.065 3166.630 541.135 ;
        RECT 0.000 537.915 3165.950 539.065 ;
        RECT 0.000 533.085 3166.630 537.915 ;
        RECT 0.000 531.935 3165.950 533.085 ;
        RECT 0.000 529.865 3166.630 531.935 ;
        RECT 0.000 528.715 3165.950 529.865 ;
        RECT 0.000 520.665 3166.630 528.715 ;
        RECT 0.000 519.515 3165.950 520.665 ;
        RECT 0.000 390.745 3166.630 519.515 ;
        RECT 0.000 389.635 3165.950 390.745 ;
        RECT 0.000 381.290 3166.630 389.635 ;
        RECT 0.000 380.735 3166.640 381.290 ;
        RECT 0.000 379.625 3165.950 380.735 ;
        RECT 3166.340 380.610 3166.640 380.735 ;
        RECT 3166.030 380.335 3166.640 380.610 ;
        RECT 0.000 368.265 3166.630 379.625 ;
        RECT 0.000 367.115 3165.950 368.265 ;
        RECT 0.000 365.505 3166.630 367.115 ;
        RECT 0.000 364.355 3165.950 365.505 ;
        RECT 0.000 362.285 3166.630 364.355 ;
        RECT 0.000 361.135 3165.950 362.285 ;
        RECT 3166.030 361.270 3166.640 361.535 ;
        RECT 3166.340 361.135 3166.640 361.270 ;
        RECT 0.000 360.590 3166.640 361.135 ;
        RECT 0.000 359.065 3166.630 360.590 ;
        RECT 0.000 357.915 3165.950 359.065 ;
        RECT 0.000 349.865 3166.630 357.915 ;
        RECT 0.000 348.715 3165.950 349.865 ;
        RECT 0.000 347.105 3166.630 348.715 ;
        RECT 0.000 345.955 3165.950 347.105 ;
        RECT 0.000 343.885 3166.630 345.955 ;
        RECT 0.000 342.735 3165.950 343.885 ;
        RECT 3166.030 342.910 3166.640 343.135 ;
        RECT 3166.340 342.735 3166.640 342.910 ;
        RECT 0.000 340.870 3166.640 342.735 ;
        RECT 0.000 340.665 3166.630 340.870 ;
        RECT 0.000 339.515 3165.950 340.665 ;
        RECT 0.000 328.245 3166.630 339.515 ;
        RECT 0.000 327.095 3165.950 328.245 ;
        RECT 0.000 325.485 3166.630 327.095 ;
        RECT 0.000 324.335 3165.950 325.485 ;
        RECT 0.000 322.265 3166.630 324.335 ;
        RECT 0.000 321.115 3165.950 322.265 ;
        RECT 0.000 319.045 3166.630 321.115 ;
        RECT 0.000 317.895 3165.950 319.045 ;
        RECT 0.000 316.285 3166.630 317.895 ;
        RECT 0.000 315.135 3165.950 316.285 ;
        RECT 0.000 313.065 3166.630 315.135 ;
        RECT 0.000 311.915 3165.950 313.065 ;
        RECT 0.000 307.085 3166.630 311.915 ;
        RECT 0.000 305.935 3165.950 307.085 ;
        RECT 0.000 303.865 3166.630 305.935 ;
        RECT 0.000 302.715 3165.950 303.865 ;
        RECT 0.000 294.665 3166.630 302.715 ;
        RECT 0.000 293.515 3165.950 294.665 ;
        RECT 0.000 268.725 3166.630 293.515 ;
        RECT 0.680 265.335 3166.630 268.725 ;
        RECT 0.000 40.635 3166.630 265.335 ;
      LAYER met4 ;
        RECT 558.970 3447.590 574.850 3478.080 ;
        RECT 582.050 3447.590 584.450 3478.080 ;
        RECT 591.650 3447.590 614.850 3478.080 ;
        RECT 622.050 3447.590 624.450 3478.080 ;
        RECT 631.650 3447.590 654.850 3478.080 ;
        RECT 662.050 3447.590 664.450 3478.080 ;
        RECT 671.650 3447.590 694.850 3478.080 ;
        RECT 702.050 3447.590 704.450 3478.080 ;
        RECT 711.650 3447.590 734.850 3478.080 ;
        RECT 742.050 3447.590 744.450 3478.080 ;
        RECT 751.650 3447.590 774.850 3478.080 ;
        RECT 782.050 3447.590 784.450 3478.080 ;
        RECT 791.650 3447.590 814.850 3478.080 ;
        RECT 822.050 3447.590 824.450 3478.080 ;
        RECT 831.650 3447.590 854.850 3478.080 ;
        RECT 862.050 3447.590 864.450 3478.080 ;
        RECT 871.650 3447.590 894.850 3478.080 ;
        RECT 902.050 3447.590 904.450 3478.080 ;
        RECT 911.650 3447.590 934.850 3478.080 ;
        RECT 942.050 3447.590 944.450 3478.080 ;
        RECT 951.650 3447.590 974.850 3478.080 ;
        RECT 982.050 3447.590 984.450 3478.080 ;
        RECT 991.650 3447.590 1014.850 3478.080 ;
        RECT 1022.050 3447.590 1024.450 3478.080 ;
        RECT 1031.650 3447.590 1054.850 3478.080 ;
        RECT 1062.050 3447.590 1064.450 3478.080 ;
        RECT 1071.650 3447.590 1094.850 3478.080 ;
        RECT 1102.050 3447.590 1104.450 3478.080 ;
        RECT 1111.650 3447.590 1134.850 3478.080 ;
        RECT 1142.050 3447.590 1144.450 3478.080 ;
        RECT 1151.650 3447.590 1174.850 3478.080 ;
        RECT 1182.050 3447.590 1184.450 3478.080 ;
        RECT 1191.650 3447.590 1214.850 3478.080 ;
        RECT 1222.050 3447.590 1224.450 3478.080 ;
        RECT 1231.650 3447.590 1254.850 3478.080 ;
        RECT 1262.050 3447.590 1264.450 3478.080 ;
        RECT 1271.650 3447.590 1294.850 3478.080 ;
        RECT 1302.050 3447.590 1304.450 3478.080 ;
        RECT 1311.650 3447.590 1334.850 3478.080 ;
        RECT 1342.050 3447.590 1344.450 3478.080 ;
        RECT 1351.650 3447.590 1374.850 3478.080 ;
        RECT 1382.050 3447.590 1384.450 3478.080 ;
        RECT 1391.650 3447.590 1414.850 3478.080 ;
        RECT 1422.050 3447.590 1424.450 3478.080 ;
        RECT 1431.650 3447.590 1454.850 3478.080 ;
        RECT 1462.050 3447.590 1464.450 3478.080 ;
        RECT 1471.650 3447.590 1494.850 3478.080 ;
        RECT 1502.050 3447.590 1504.450 3478.080 ;
        RECT 1511.650 3447.590 1534.850 3478.080 ;
        RECT 1542.050 3447.590 1544.450 3478.080 ;
        RECT 1551.650 3447.590 1574.850 3478.080 ;
        RECT 1582.050 3447.590 1584.450 3478.080 ;
        RECT 1591.650 3447.590 1614.850 3478.080 ;
        RECT 1622.050 3447.590 1624.450 3478.080 ;
        RECT 1631.650 3447.590 1654.850 3478.080 ;
        RECT 1662.050 3447.590 1664.450 3478.080 ;
        RECT 1671.650 3447.590 1694.850 3478.080 ;
        RECT 1702.050 3447.590 1704.450 3478.080 ;
        RECT 1711.650 3447.590 1734.850 3478.080 ;
        RECT 1742.050 3447.590 1744.450 3478.080 ;
        RECT 1751.650 3447.590 1774.850 3478.080 ;
        RECT 1782.050 3447.590 1784.450 3478.080 ;
        RECT 1791.650 3447.590 1814.850 3478.080 ;
        RECT 1822.050 3447.590 1824.450 3478.080 ;
        RECT 1831.650 3447.590 1854.850 3478.080 ;
        RECT 1862.050 3447.590 1864.450 3478.080 ;
        RECT 1871.650 3447.590 1894.850 3478.080 ;
        RECT 1902.050 3447.590 1904.450 3478.080 ;
        RECT 1911.650 3447.590 1934.850 3478.080 ;
        RECT 1942.050 3447.590 1944.450 3478.080 ;
        RECT 1951.650 3447.590 1974.850 3478.080 ;
        RECT 1982.050 3447.590 1984.450 3478.080 ;
        RECT 1991.650 3447.590 2014.850 3478.080 ;
        RECT 2022.050 3447.590 2024.450 3478.080 ;
        RECT 2031.650 3447.590 2054.850 3478.080 ;
        RECT 2062.050 3447.590 2064.450 3478.080 ;
        RECT 2071.650 3447.590 2094.850 3478.080 ;
        RECT 2102.050 3447.590 2104.450 3478.080 ;
        RECT 2111.650 3447.590 2134.850 3478.080 ;
        RECT 2142.050 3447.590 2144.450 3478.080 ;
        RECT 2151.650 3447.590 2174.850 3478.080 ;
        RECT 2182.050 3447.590 2184.450 3478.080 ;
        RECT 2191.650 3447.590 2214.850 3478.080 ;
        RECT 2222.050 3447.590 2224.450 3478.080 ;
        RECT 2231.650 3447.590 2254.850 3478.080 ;
        RECT 2262.050 3447.590 2264.450 3478.080 ;
        RECT 2271.650 3447.590 2294.850 3478.080 ;
        RECT 2302.050 3447.590 2304.450 3478.080 ;
        RECT 2311.650 3447.590 2334.850 3478.080 ;
        RECT 2342.050 3447.590 2344.450 3478.080 ;
        RECT 2351.650 3447.590 2374.850 3478.080 ;
        RECT 2382.050 3447.590 2384.450 3478.080 ;
        RECT 2391.650 3447.590 2414.850 3478.080 ;
        RECT 2422.050 3447.590 2424.450 3478.080 ;
        RECT 2431.650 3447.590 2454.850 3478.080 ;
        RECT 2462.050 3447.590 2464.450 3478.080 ;
        RECT 2471.650 3447.590 2494.850 3478.080 ;
        RECT 2502.050 3447.590 2504.450 3478.080 ;
        RECT 2511.650 3447.590 2534.850 3478.080 ;
        RECT 2542.050 3447.590 2544.450 3478.080 ;
        RECT 2551.650 3447.590 2574.850 3478.080 ;
        RECT 2582.050 3447.590 2584.450 3478.080 ;
        RECT 2591.650 3447.590 2614.850 3478.080 ;
        RECT 2622.050 3447.590 2624.450 3478.080 ;
        RECT 2631.650 3447.590 2654.850 3478.080 ;
        RECT 2662.050 3447.590 2664.450 3478.080 ;
        RECT 2671.650 3447.590 2694.850 3478.080 ;
        RECT 2702.050 3447.590 2704.450 3478.080 ;
        RECT 2711.650 3447.590 2734.850 3478.080 ;
        RECT 558.970 2051.275 2736.545 3447.590 ;
        RECT 558.970 2000.640 574.850 2051.275 ;
        RECT 582.050 2000.640 584.450 2051.275 ;
        RECT 591.650 2000.640 614.850 2051.275 ;
        RECT 622.050 2000.640 624.450 2051.275 ;
        RECT 631.650 2000.640 654.850 2051.275 ;
        RECT 662.050 2000.640 664.450 2051.275 ;
        RECT 671.650 2000.640 694.850 2051.275 ;
        RECT 702.050 2000.640 704.450 2051.275 ;
        RECT 711.650 2000.640 734.850 2051.275 ;
        RECT 742.050 2000.640 744.450 2051.275 ;
        RECT 751.650 2000.640 774.850 2051.275 ;
        RECT 782.050 2000.640 784.450 2051.275 ;
        RECT 791.650 2000.640 814.850 2051.275 ;
        RECT 822.050 2000.640 824.450 2051.275 ;
        RECT 831.650 2000.640 854.850 2051.275 ;
        RECT 862.050 2000.640 864.450 2051.275 ;
        RECT 871.650 2000.640 894.850 2051.275 ;
        RECT 902.050 2000.640 904.450 2051.275 ;
        RECT 911.650 2000.640 934.850 2051.275 ;
        RECT 942.050 2000.640 944.450 2051.275 ;
        RECT 951.650 2000.640 974.850 2051.275 ;
        RECT 982.050 2000.640 984.450 2051.275 ;
        RECT 991.650 2000.640 1014.850 2051.275 ;
        RECT 1022.050 2000.640 1024.450 2051.275 ;
        RECT 1031.650 2000.640 1054.850 2051.275 ;
        RECT 1062.050 2000.640 1064.450 2051.275 ;
        RECT 1071.650 2000.640 1094.850 2051.275 ;
        RECT 1102.050 2000.640 1104.450 2051.275 ;
        RECT 1111.650 2000.640 1134.850 2051.275 ;
        RECT 1142.050 2000.640 1144.450 2051.275 ;
        RECT 1151.650 2000.640 1174.850 2051.275 ;
        RECT 1182.050 2000.640 1184.450 2051.275 ;
        RECT 1191.650 2000.640 1214.850 2051.275 ;
        RECT 1222.050 2000.640 1224.450 2051.275 ;
        RECT 1231.650 2000.640 1254.850 2051.275 ;
        RECT 1262.050 2000.640 1264.450 2051.275 ;
        RECT 1271.650 2000.640 1294.850 2051.275 ;
        RECT 1302.050 2000.640 1304.450 2051.275 ;
        RECT 1311.650 2000.640 1334.850 2051.275 ;
        RECT 1342.050 2000.640 1344.450 2051.275 ;
        RECT 1351.650 2000.640 1374.850 2051.275 ;
        RECT 1382.050 2000.640 1384.450 2051.275 ;
        RECT 1391.650 2000.640 1414.850 2051.275 ;
        RECT 1422.050 2000.640 1424.450 2051.275 ;
        RECT 1431.650 2000.640 1454.850 2051.275 ;
        RECT 1462.050 2000.640 1464.450 2051.275 ;
        RECT 1471.650 2000.640 1494.850 2051.275 ;
        RECT 1502.050 2000.640 1504.450 2051.275 ;
        RECT 1511.650 2000.640 1534.850 2051.275 ;
        RECT 1542.050 2000.640 1544.450 2051.275 ;
        RECT 1551.650 2000.640 1574.850 2051.275 ;
        RECT 1582.050 2000.640 1584.450 2051.275 ;
        RECT 1591.650 2000.640 1614.850 2051.275 ;
        RECT 1622.050 2000.640 1624.450 2051.275 ;
        RECT 1631.650 2000.640 1654.850 2051.275 ;
        RECT 1662.050 2000.640 1664.450 2051.275 ;
        RECT 1671.650 2000.640 1694.850 2051.275 ;
        RECT 1702.050 2000.640 1704.450 2051.275 ;
        RECT 1711.650 2000.640 1734.850 2051.275 ;
        RECT 1742.050 2000.640 1744.450 2051.275 ;
        RECT 1751.650 2000.640 1774.850 2051.275 ;
        RECT 1782.050 2000.640 1784.450 2051.275 ;
        RECT 1791.650 2000.640 1814.850 2051.275 ;
        RECT 1822.050 2000.640 1824.450 2051.275 ;
        RECT 1831.650 2000.640 1854.850 2051.275 ;
        RECT 1862.050 2000.640 1864.450 2051.275 ;
        RECT 1871.650 2000.640 1894.850 2051.275 ;
        RECT 1902.050 2000.640 1904.450 2051.275 ;
        RECT 1911.650 2000.640 1934.850 2051.275 ;
        RECT 1942.050 2000.640 1944.450 2051.275 ;
        RECT 1951.650 2000.640 1974.850 2051.275 ;
        RECT 1982.050 2000.640 1984.450 2051.275 ;
        RECT 1991.650 2000.640 2014.850 2051.275 ;
        RECT 2022.050 2000.640 2024.450 2051.275 ;
        RECT 2031.650 2000.640 2054.850 2051.275 ;
        RECT 2062.050 2000.640 2064.450 2051.275 ;
        RECT 2071.650 2000.640 2094.850 2051.275 ;
        RECT 2102.050 2000.640 2104.450 2051.275 ;
        RECT 2111.650 2000.640 2134.850 2051.275 ;
        RECT 2142.050 2000.640 2144.450 2051.275 ;
        RECT 2151.650 2000.640 2174.850 2051.275 ;
        RECT 2182.050 2000.640 2184.450 2051.275 ;
        RECT 2191.650 2000.640 2214.850 2051.275 ;
        RECT 2222.050 2000.640 2224.450 2051.275 ;
        RECT 2231.650 2000.640 2254.850 2051.275 ;
        RECT 2262.050 2000.640 2264.450 2051.275 ;
        RECT 2271.650 2000.640 2294.850 2051.275 ;
        RECT 2302.050 2000.640 2304.450 2051.275 ;
        RECT 2311.650 2000.640 2334.850 2051.275 ;
        RECT 2342.050 2000.640 2344.450 2051.275 ;
        RECT 2351.650 2000.640 2374.850 2051.275 ;
        RECT 2382.050 2000.640 2384.450 2051.275 ;
        RECT 2391.650 2000.640 2414.850 2051.275 ;
        RECT 2422.050 2000.640 2424.450 2051.275 ;
        RECT 2431.650 2000.640 2454.850 2051.275 ;
        RECT 2462.050 2000.640 2464.450 2051.275 ;
        RECT 2471.650 2000.640 2494.850 2051.275 ;
        RECT 2502.050 2000.640 2504.450 2051.275 ;
        RECT 2511.650 2000.640 2534.850 2051.275 ;
        RECT 2542.050 2000.640 2544.450 2051.275 ;
        RECT 2551.650 2000.640 2574.850 2051.275 ;
        RECT 2582.050 2000.640 2584.450 2051.275 ;
        RECT 2591.650 2000.640 2614.850 2051.275 ;
        RECT 2622.050 2000.640 2624.450 2051.275 ;
        RECT 2631.650 2000.640 2654.850 2051.275 ;
        RECT 2662.050 2000.640 2664.450 2051.275 ;
        RECT 2671.650 2000.640 2694.850 2051.275 ;
        RECT 2702.050 2000.640 2704.450 2051.275 ;
        RECT 2711.650 2000.640 2734.850 2051.275 ;
      LAYER met5 ;
        RECT 555.280 3438.030 2744.440 3452.530 ;
        RECT 625.460 3418.830 2404.700 3438.030 ;
        RECT 555.280 3398.030 2744.440 3418.830 ;
        RECT 625.460 3378.830 2404.700 3398.030 ;
        RECT 555.280 3358.030 2744.440 3378.830 ;
        RECT 625.460 3338.830 2404.700 3358.030 ;
        RECT 555.280 3318.030 2744.440 3338.830 ;
        RECT 625.460 3298.830 2404.700 3318.030 ;
        RECT 555.280 3278.030 2744.440 3298.830 ;
        RECT 625.460 3258.830 2404.700 3278.030 ;
        RECT 555.280 3238.030 2744.440 3258.830 ;
        RECT 625.460 3218.830 2404.700 3238.030 ;
        RECT 555.280 3198.030 2744.440 3218.830 ;
        RECT 625.460 3178.830 2404.700 3198.030 ;
        RECT 555.280 3158.030 2744.440 3178.830 ;
        RECT 625.460 3138.830 2404.700 3158.030 ;
        RECT 555.280 3118.030 2744.440 3138.830 ;
        RECT 625.460 3098.830 2404.700 3118.030 ;
        RECT 555.280 3078.030 2744.440 3098.830 ;
        RECT 625.460 3058.830 2404.700 3078.030 ;
        RECT 555.280 3038.030 2744.440 3058.830 ;
        RECT 625.460 3018.830 2404.700 3038.030 ;
        RECT 555.280 2998.030 2744.440 3018.830 ;
        RECT 625.460 2978.830 2404.700 2998.030 ;
        RECT 555.280 2958.030 2744.440 2978.830 ;
        RECT 625.460 2938.830 2404.700 2958.030 ;
        RECT 555.280 2918.030 2744.440 2938.830 ;
        RECT 625.460 2898.830 2404.700 2918.030 ;
        RECT 555.280 2878.030 2744.440 2898.830 ;
        RECT 625.460 2858.830 2404.700 2878.030 ;
        RECT 555.280 2838.030 2744.440 2858.830 ;
        RECT 625.460 2818.830 2404.700 2838.030 ;
        RECT 555.280 2798.030 2744.440 2818.830 ;
        RECT 625.460 2778.830 2404.700 2798.030 ;
        RECT 555.280 2758.030 2744.440 2778.830 ;
        RECT 625.460 2738.830 2404.700 2758.030 ;
        RECT 555.280 2718.030 2744.440 2738.830 ;
        RECT 625.460 2698.830 2404.700 2718.030 ;
        RECT 555.280 2678.030 2744.440 2698.830 ;
        RECT 625.460 2658.830 2404.700 2678.030 ;
        RECT 555.280 2638.030 2744.440 2658.830 ;
        RECT 625.460 2618.830 2404.700 2638.030 ;
        RECT 555.280 2598.030 2744.440 2618.830 ;
        RECT 625.460 2578.830 2404.700 2598.030 ;
        RECT 555.280 2558.030 2744.440 2578.830 ;
        RECT 625.460 2538.830 2404.700 2558.030 ;
        RECT 555.280 2518.030 2744.440 2538.830 ;
        RECT 625.460 2498.830 2404.700 2518.030 ;
        RECT 555.280 2478.030 2744.440 2498.830 ;
        RECT 555.280 2438.030 2744.440 2458.830 ;
        RECT 555.280 2398.030 2744.440 2418.830 ;
        RECT 555.280 2358.030 2744.440 2378.830 ;
        RECT 555.280 2318.030 2744.440 2338.830 ;
        RECT 555.280 2278.030 2744.440 2298.830 ;
        RECT 555.280 2238.030 2744.440 2258.830 ;
        RECT 555.280 2198.030 2744.440 2218.830 ;
        RECT 555.280 2158.030 2744.440 2178.830 ;
        RECT 555.280 2118.030 2744.440 2138.830 ;
        RECT 555.280 2078.030 2744.440 2098.830 ;
        RECT 555.280 2038.030 2744.440 2058.830 ;
        RECT 555.280 2004.330 2744.440 2018.830 ;
  END
END openframe_project_wrapper
END LIBRARY

