magic
tech sky130A
magscale 1 2
timestamp 1685898580
<< obsli1 >>
rect 1104 2159 438840 277457
<< obsm1 >>
rect 14 1776 438840 277704
<< metal2 >>
rect 3330 279520 3386 280000
rect 7378 279520 7434 280000
rect 11426 279520 11482 280000
rect 15474 279520 15530 280000
rect 19522 279520 19578 280000
rect 23570 279520 23626 280000
rect 27618 279520 27674 280000
rect 31666 279520 31722 280000
rect 35714 279520 35770 280000
rect 39762 279520 39818 280000
rect 43810 279520 43866 280000
rect 47858 279520 47914 280000
rect 51906 279520 51962 280000
rect 55954 279520 56010 280000
rect 60002 279520 60058 280000
rect 64050 279520 64106 280000
rect 68098 279520 68154 280000
rect 72146 279520 72202 280000
rect 76194 279520 76250 280000
rect 80242 279520 80298 280000
rect 84290 279520 84346 280000
rect 88338 279520 88394 280000
rect 92386 279520 92442 280000
rect 96434 279520 96490 280000
rect 100482 279520 100538 280000
rect 104530 279520 104586 280000
rect 108578 279520 108634 280000
rect 112626 279520 112682 280000
rect 116674 279520 116730 280000
rect 120722 279520 120778 280000
rect 124770 279520 124826 280000
rect 128818 279520 128874 280000
rect 132866 279520 132922 280000
rect 136914 279520 136970 280000
rect 140962 279520 141018 280000
rect 145010 279520 145066 280000
rect 149058 279520 149114 280000
rect 153106 279520 153162 280000
rect 157154 279520 157210 280000
rect 161202 279520 161258 280000
rect 165250 279520 165306 280000
rect 169298 279520 169354 280000
rect 173346 279520 173402 280000
rect 177394 279520 177450 280000
rect 181442 279520 181498 280000
rect 185490 279520 185546 280000
rect 189538 279520 189594 280000
rect 193586 279520 193642 280000
rect 197634 279520 197690 280000
rect 201682 279520 201738 280000
rect 205730 279520 205786 280000
rect 209778 279520 209834 280000
rect 213826 279520 213882 280000
rect 217874 279520 217930 280000
rect 221922 279520 221978 280000
rect 225970 279520 226026 280000
rect 230018 279520 230074 280000
rect 234066 279520 234122 280000
rect 238114 279520 238170 280000
rect 242162 279520 242218 280000
rect 246210 279520 246266 280000
rect 250258 279520 250314 280000
rect 254306 279520 254362 280000
rect 258354 279520 258410 280000
rect 262402 279520 262458 280000
rect 266450 279520 266506 280000
rect 270498 279520 270554 280000
rect 274546 279520 274602 280000
rect 278594 279520 278650 280000
rect 282642 279520 282698 280000
rect 286690 279520 286746 280000
rect 290738 279520 290794 280000
rect 294786 279520 294842 280000
rect 298834 279520 298890 280000
rect 302882 279520 302938 280000
rect 306930 279520 306986 280000
rect 310978 279520 311034 280000
rect 315026 279520 315082 280000
rect 319074 279520 319130 280000
rect 323122 279520 323178 280000
rect 327170 279520 327226 280000
rect 331218 279520 331274 280000
rect 335266 279520 335322 280000
rect 339314 279520 339370 280000
rect 343362 279520 343418 280000
rect 347410 279520 347466 280000
rect 351458 279520 351514 280000
rect 355506 279520 355562 280000
rect 359554 279520 359610 280000
rect 363602 279520 363658 280000
rect 367650 279520 367706 280000
rect 371698 279520 371754 280000
rect 375746 279520 375802 280000
rect 379794 279520 379850 280000
rect 383842 279520 383898 280000
rect 387890 279520 387946 280000
rect 391938 279520 391994 280000
rect 395986 279520 396042 280000
rect 400034 279520 400090 280000
rect 404082 279520 404138 280000
rect 408130 279520 408186 280000
rect 412178 279520 412234 280000
rect 416226 279520 416282 280000
rect 420274 279520 420330 280000
rect 424322 279520 424378 280000
rect 428370 279520 428426 280000
rect 432418 279520 432474 280000
rect 436466 279520 436522 280000
rect 4618 0 4674 480
rect 8758 0 8814 480
rect 12898 0 12954 480
rect 17038 0 17094 480
rect 21178 0 21234 480
rect 25318 0 25374 480
rect 29458 0 29514 480
rect 33598 0 33654 480
rect 37738 0 37794 480
rect 41878 0 41934 480
rect 46018 0 46074 480
rect 50158 0 50214 480
rect 54298 0 54354 480
rect 58438 0 58494 480
rect 62578 0 62634 480
rect 66718 0 66774 480
rect 70858 0 70914 480
rect 74998 0 75054 480
rect 79138 0 79194 480
rect 83278 0 83334 480
rect 87418 0 87474 480
rect 91558 0 91614 480
rect 95698 0 95754 480
rect 99838 0 99894 480
rect 103978 0 104034 480
rect 108118 0 108174 480
rect 112258 0 112314 480
rect 116398 0 116454 480
rect 120538 0 120594 480
rect 124678 0 124734 480
rect 128818 0 128874 480
rect 132958 0 133014 480
rect 137098 0 137154 480
rect 141238 0 141294 480
rect 145378 0 145434 480
rect 149518 0 149574 480
rect 153658 0 153714 480
rect 157798 0 157854 480
rect 161938 0 161994 480
rect 166078 0 166134 480
rect 170218 0 170274 480
rect 174358 0 174414 480
rect 178498 0 178554 480
rect 182638 0 182694 480
rect 186778 0 186834 480
rect 190918 0 190974 480
rect 195058 0 195114 480
rect 199198 0 199254 480
rect 203338 0 203394 480
rect 207478 0 207534 480
rect 211618 0 211674 480
rect 215758 0 215814 480
rect 219898 0 219954 480
rect 224038 0 224094 480
rect 228178 0 228234 480
rect 232318 0 232374 480
rect 236458 0 236514 480
rect 240598 0 240654 480
rect 244738 0 244794 480
rect 248878 0 248934 480
rect 253018 0 253074 480
rect 257158 0 257214 480
rect 261298 0 261354 480
rect 265438 0 265494 480
rect 269578 0 269634 480
rect 273718 0 273774 480
rect 277858 0 277914 480
rect 281998 0 282054 480
rect 286138 0 286194 480
rect 290278 0 290334 480
rect 294418 0 294474 480
rect 298558 0 298614 480
rect 302698 0 302754 480
rect 306838 0 306894 480
rect 310978 0 311034 480
rect 315118 0 315174 480
rect 319258 0 319314 480
rect 323398 0 323454 480
rect 327538 0 327594 480
rect 331678 0 331734 480
rect 335818 0 335874 480
rect 339958 0 340014 480
rect 344098 0 344154 480
rect 348238 0 348294 480
rect 352378 0 352434 480
rect 356518 0 356574 480
rect 360658 0 360714 480
rect 364798 0 364854 480
rect 368938 0 368994 480
rect 373078 0 373134 480
rect 377218 0 377274 480
rect 381358 0 381414 480
rect 385498 0 385554 480
rect 389638 0 389694 480
rect 393778 0 393834 480
rect 397918 0 397974 480
rect 402058 0 402114 480
rect 406198 0 406254 480
rect 410338 0 410394 480
rect 414478 0 414534 480
rect 418618 0 418674 480
rect 422758 0 422814 480
rect 426898 0 426954 480
rect 431038 0 431094 480
rect 435178 0 435234 480
<< obsm2 >>
rect 18 279464 3274 279562
rect 3442 279464 7322 279562
rect 7490 279464 11370 279562
rect 11538 279464 15418 279562
rect 15586 279464 19466 279562
rect 19634 279464 23514 279562
rect 23682 279464 27562 279562
rect 27730 279464 31610 279562
rect 31778 279464 35658 279562
rect 35826 279464 39706 279562
rect 39874 279464 43754 279562
rect 43922 279464 47802 279562
rect 47970 279464 51850 279562
rect 52018 279464 55898 279562
rect 56066 279464 59946 279562
rect 60114 279464 63994 279562
rect 64162 279464 68042 279562
rect 68210 279464 72090 279562
rect 72258 279464 76138 279562
rect 76306 279464 80186 279562
rect 80354 279464 84234 279562
rect 84402 279464 88282 279562
rect 88450 279464 92330 279562
rect 92498 279464 96378 279562
rect 96546 279464 100426 279562
rect 100594 279464 104474 279562
rect 104642 279464 108522 279562
rect 108690 279464 112570 279562
rect 112738 279464 116618 279562
rect 116786 279464 120666 279562
rect 120834 279464 124714 279562
rect 124882 279464 128762 279562
rect 128930 279464 132810 279562
rect 132978 279464 136858 279562
rect 137026 279464 140906 279562
rect 141074 279464 144954 279562
rect 145122 279464 149002 279562
rect 149170 279464 153050 279562
rect 153218 279464 157098 279562
rect 157266 279464 161146 279562
rect 161314 279464 165194 279562
rect 165362 279464 169242 279562
rect 169410 279464 173290 279562
rect 173458 279464 177338 279562
rect 177506 279464 181386 279562
rect 181554 279464 185434 279562
rect 185602 279464 189482 279562
rect 189650 279464 193530 279562
rect 193698 279464 197578 279562
rect 197746 279464 201626 279562
rect 201794 279464 205674 279562
rect 205842 279464 209722 279562
rect 209890 279464 213770 279562
rect 213938 279464 217818 279562
rect 217986 279464 221866 279562
rect 222034 279464 225914 279562
rect 226082 279464 229962 279562
rect 230130 279464 234010 279562
rect 234178 279464 238058 279562
rect 238226 279464 242106 279562
rect 242274 279464 246154 279562
rect 246322 279464 250202 279562
rect 250370 279464 254250 279562
rect 254418 279464 258298 279562
rect 258466 279464 262346 279562
rect 262514 279464 266394 279562
rect 266562 279464 270442 279562
rect 270610 279464 274490 279562
rect 274658 279464 278538 279562
rect 278706 279464 282586 279562
rect 282754 279464 286634 279562
rect 286802 279464 290682 279562
rect 290850 279464 294730 279562
rect 294898 279464 298778 279562
rect 298946 279464 302826 279562
rect 302994 279464 306874 279562
rect 307042 279464 310922 279562
rect 311090 279464 314970 279562
rect 315138 279464 319018 279562
rect 319186 279464 323066 279562
rect 323234 279464 327114 279562
rect 327282 279464 331162 279562
rect 331330 279464 335210 279562
rect 335378 279464 339258 279562
rect 339426 279464 343306 279562
rect 343474 279464 347354 279562
rect 347522 279464 351402 279562
rect 351570 279464 355450 279562
rect 355618 279464 359498 279562
rect 359666 279464 363546 279562
rect 363714 279464 367594 279562
rect 367762 279464 371642 279562
rect 371810 279464 375690 279562
rect 375858 279464 379738 279562
rect 379906 279464 383786 279562
rect 383954 279464 387834 279562
rect 388002 279464 391882 279562
rect 392050 279464 395930 279562
rect 396098 279464 399978 279562
rect 400146 279464 404026 279562
rect 404194 279464 408074 279562
rect 408242 279464 412122 279562
rect 412290 279464 416170 279562
rect 416338 279464 420218 279562
rect 420386 279464 424266 279562
rect 424434 279464 428314 279562
rect 428482 279464 432362 279562
rect 432530 279464 436410 279562
rect 436578 279464 438822 279562
rect 18 536 438822 279464
rect 18 326 4562 536
rect 4730 326 8702 536
rect 8870 326 12842 536
rect 13010 326 16982 536
rect 17150 326 21122 536
rect 21290 326 25262 536
rect 25430 326 29402 536
rect 29570 326 33542 536
rect 33710 326 37682 536
rect 37850 326 41822 536
rect 41990 326 45962 536
rect 46130 326 50102 536
rect 50270 326 54242 536
rect 54410 326 58382 536
rect 58550 326 62522 536
rect 62690 326 66662 536
rect 66830 326 70802 536
rect 70970 326 74942 536
rect 75110 326 79082 536
rect 79250 326 83222 536
rect 83390 326 87362 536
rect 87530 326 91502 536
rect 91670 326 95642 536
rect 95810 326 99782 536
rect 99950 326 103922 536
rect 104090 326 108062 536
rect 108230 326 112202 536
rect 112370 326 116342 536
rect 116510 326 120482 536
rect 120650 326 124622 536
rect 124790 326 128762 536
rect 128930 326 132902 536
rect 133070 326 137042 536
rect 137210 326 141182 536
rect 141350 326 145322 536
rect 145490 326 149462 536
rect 149630 326 153602 536
rect 153770 326 157742 536
rect 157910 326 161882 536
rect 162050 326 166022 536
rect 166190 326 170162 536
rect 170330 326 174302 536
rect 174470 326 178442 536
rect 178610 326 182582 536
rect 182750 326 186722 536
rect 186890 326 190862 536
rect 191030 326 195002 536
rect 195170 326 199142 536
rect 199310 326 203282 536
rect 203450 326 207422 536
rect 207590 326 211562 536
rect 211730 326 215702 536
rect 215870 326 219842 536
rect 220010 326 223982 536
rect 224150 326 228122 536
rect 228290 326 232262 536
rect 232430 326 236402 536
rect 236570 326 240542 536
rect 240710 326 244682 536
rect 244850 326 248822 536
rect 248990 326 252962 536
rect 253130 326 257102 536
rect 257270 326 261242 536
rect 261410 326 265382 536
rect 265550 326 269522 536
rect 269690 326 273662 536
rect 273830 326 277802 536
rect 277970 326 281942 536
rect 282110 326 286082 536
rect 286250 326 290222 536
rect 290390 326 294362 536
rect 294530 326 298502 536
rect 298670 326 302642 536
rect 302810 326 306782 536
rect 306950 326 310922 536
rect 311090 326 315062 536
rect 315230 326 319202 536
rect 319370 326 323342 536
rect 323510 326 327482 536
rect 327650 326 331622 536
rect 331790 326 335762 536
rect 335930 326 339902 536
rect 340070 326 344042 536
rect 344210 326 348182 536
rect 348350 326 352322 536
rect 352490 326 356462 536
rect 356630 326 360602 536
rect 360770 326 364742 536
rect 364910 326 368882 536
rect 369050 326 373022 536
rect 373190 326 377162 536
rect 377330 326 381302 536
rect 381470 326 385442 536
rect 385610 326 389582 536
rect 389750 326 393722 536
rect 393890 326 397862 536
rect 398030 326 402002 536
rect 402170 326 406142 536
rect 406310 326 410282 536
rect 410450 326 414422 536
rect 414590 326 418562 536
rect 418730 326 422702 536
rect 422870 326 426842 536
rect 427010 326 430982 536
rect 431150 326 435122 536
rect 435290 326 438822 536
<< metal3 >>
rect 0 277720 480 277840
rect 0 276088 480 276208
rect 0 274456 480 274576
rect 0 272824 480 272944
rect 0 271192 480 271312
rect 0 269560 480 269680
rect 0 267928 480 268048
rect 0 266296 480 266416
rect 0 264664 480 264784
rect 0 263032 480 263152
rect 439520 261672 440000 261792
rect 0 261400 480 261520
rect 439520 260312 440000 260432
rect 0 259768 480 259888
rect 439520 258952 440000 259072
rect 0 258136 480 258256
rect 439520 257592 440000 257712
rect 0 256504 480 256624
rect 439520 256232 440000 256352
rect 0 254872 480 254992
rect 439520 254872 440000 254992
rect 439520 253512 440000 253632
rect 0 253240 480 253360
rect 439520 252152 440000 252272
rect 0 251608 480 251728
rect 439520 250792 440000 250912
rect 0 249976 480 250096
rect 439520 249432 440000 249552
rect 0 248344 480 248464
rect 439520 248072 440000 248192
rect 0 246712 480 246832
rect 439520 246712 440000 246832
rect 439520 245352 440000 245472
rect 0 245080 480 245200
rect 439520 243992 440000 244112
rect 0 243448 480 243568
rect 439520 242632 440000 242752
rect 0 241816 480 241936
rect 439520 241272 440000 241392
rect 0 240184 480 240304
rect 439520 239912 440000 240032
rect 0 238552 480 238672
rect 439520 238552 440000 238672
rect 439520 237192 440000 237312
rect 0 236920 480 237040
rect 439520 235832 440000 235952
rect 0 235288 480 235408
rect 439520 234472 440000 234592
rect 0 233656 480 233776
rect 439520 233112 440000 233232
rect 0 232024 480 232144
rect 439520 231752 440000 231872
rect 0 230392 480 230512
rect 439520 230392 440000 230512
rect 439520 229032 440000 229152
rect 0 228760 480 228880
rect 439520 227672 440000 227792
rect 0 227128 480 227248
rect 439520 226312 440000 226432
rect 0 225496 480 225616
rect 439520 224952 440000 225072
rect 0 223864 480 223984
rect 439520 223592 440000 223712
rect 0 222232 480 222352
rect 439520 222232 440000 222352
rect 439520 220872 440000 220992
rect 0 220600 480 220720
rect 439520 219512 440000 219632
rect 0 218968 480 219088
rect 439520 218152 440000 218272
rect 0 217336 480 217456
rect 439520 216792 440000 216912
rect 0 215704 480 215824
rect 439520 215432 440000 215552
rect 0 214072 480 214192
rect 439520 214072 440000 214192
rect 439520 212712 440000 212832
rect 0 212440 480 212560
rect 439520 211352 440000 211472
rect 0 210808 480 210928
rect 439520 209992 440000 210112
rect 0 209176 480 209296
rect 439520 208632 440000 208752
rect 0 207544 480 207664
rect 439520 207272 440000 207392
rect 0 205912 480 206032
rect 439520 205912 440000 206032
rect 439520 204552 440000 204672
rect 0 204280 480 204400
rect 439520 203192 440000 203312
rect 0 202648 480 202768
rect 439520 201832 440000 201952
rect 0 201016 480 201136
rect 439520 200472 440000 200592
rect 0 199384 480 199504
rect 439520 199112 440000 199232
rect 0 197752 480 197872
rect 439520 197752 440000 197872
rect 439520 196392 440000 196512
rect 0 196120 480 196240
rect 439520 195032 440000 195152
rect 0 194488 480 194608
rect 439520 193672 440000 193792
rect 0 192856 480 192976
rect 439520 192312 440000 192432
rect 0 191224 480 191344
rect 439520 190952 440000 191072
rect 0 189592 480 189712
rect 439520 189592 440000 189712
rect 439520 188232 440000 188352
rect 0 187960 480 188080
rect 439520 186872 440000 186992
rect 0 186328 480 186448
rect 439520 185512 440000 185632
rect 0 184696 480 184816
rect 439520 184152 440000 184272
rect 0 183064 480 183184
rect 439520 182792 440000 182912
rect 0 181432 480 181552
rect 439520 181432 440000 181552
rect 439520 180072 440000 180192
rect 0 179800 480 179920
rect 439520 178712 440000 178832
rect 0 178168 480 178288
rect 439520 177352 440000 177472
rect 0 176536 480 176656
rect 439520 175992 440000 176112
rect 0 174904 480 175024
rect 439520 174632 440000 174752
rect 0 173272 480 173392
rect 439520 173272 440000 173392
rect 439520 171912 440000 172032
rect 0 171640 480 171760
rect 439520 170552 440000 170672
rect 0 170008 480 170128
rect 439520 169192 440000 169312
rect 0 168376 480 168496
rect 439520 167832 440000 167952
rect 0 166744 480 166864
rect 439520 166472 440000 166592
rect 0 165112 480 165232
rect 439520 165112 440000 165232
rect 439520 163752 440000 163872
rect 0 163480 480 163600
rect 439520 162392 440000 162512
rect 0 161848 480 161968
rect 439520 161032 440000 161152
rect 0 160216 480 160336
rect 439520 159672 440000 159792
rect 0 158584 480 158704
rect 439520 158312 440000 158432
rect 0 156952 480 157072
rect 439520 156952 440000 157072
rect 439520 155592 440000 155712
rect 0 155320 480 155440
rect 439520 154232 440000 154352
rect 0 153688 480 153808
rect 439520 152872 440000 152992
rect 0 152056 480 152176
rect 439520 151512 440000 151632
rect 0 150424 480 150544
rect 439520 150152 440000 150272
rect 0 148792 480 148912
rect 439520 148792 440000 148912
rect 439520 147432 440000 147552
rect 0 147160 480 147280
rect 439520 146072 440000 146192
rect 0 145528 480 145648
rect 439520 144712 440000 144832
rect 0 143896 480 144016
rect 439520 143352 440000 143472
rect 0 142264 480 142384
rect 439520 141992 440000 142112
rect 0 140632 480 140752
rect 439520 140632 440000 140752
rect 439520 139272 440000 139392
rect 0 139000 480 139120
rect 439520 137912 440000 138032
rect 0 137368 480 137488
rect 439520 136552 440000 136672
rect 0 135736 480 135856
rect 439520 135192 440000 135312
rect 0 134104 480 134224
rect 439520 133832 440000 133952
rect 0 132472 480 132592
rect 439520 132472 440000 132592
rect 439520 131112 440000 131232
rect 0 130840 480 130960
rect 439520 129752 440000 129872
rect 0 129208 480 129328
rect 439520 128392 440000 128512
rect 0 127576 480 127696
rect 439520 127032 440000 127152
rect 0 125944 480 126064
rect 439520 125672 440000 125792
rect 0 124312 480 124432
rect 439520 124312 440000 124432
rect 439520 122952 440000 123072
rect 0 122680 480 122800
rect 439520 121592 440000 121712
rect 0 121048 480 121168
rect 439520 120232 440000 120352
rect 0 119416 480 119536
rect 439520 118872 440000 118992
rect 0 117784 480 117904
rect 439520 117512 440000 117632
rect 0 116152 480 116272
rect 439520 116152 440000 116272
rect 439520 114792 440000 114912
rect 0 114520 480 114640
rect 439520 113432 440000 113552
rect 0 112888 480 113008
rect 439520 112072 440000 112192
rect 0 111256 480 111376
rect 439520 110712 440000 110832
rect 0 109624 480 109744
rect 439520 109352 440000 109472
rect 0 107992 480 108112
rect 439520 107992 440000 108112
rect 439520 106632 440000 106752
rect 0 106360 480 106480
rect 439520 105272 440000 105392
rect 0 104728 480 104848
rect 439520 103912 440000 104032
rect 0 103096 480 103216
rect 439520 102552 440000 102672
rect 0 101464 480 101584
rect 439520 101192 440000 101312
rect 0 99832 480 99952
rect 439520 99832 440000 99952
rect 439520 98472 440000 98592
rect 0 98200 480 98320
rect 439520 97112 440000 97232
rect 0 96568 480 96688
rect 439520 95752 440000 95872
rect 0 94936 480 95056
rect 439520 94392 440000 94512
rect 0 93304 480 93424
rect 439520 93032 440000 93152
rect 0 91672 480 91792
rect 439520 91672 440000 91792
rect 439520 90312 440000 90432
rect 0 90040 480 90160
rect 439520 88952 440000 89072
rect 0 88408 480 88528
rect 439520 87592 440000 87712
rect 0 86776 480 86896
rect 439520 86232 440000 86352
rect 0 85144 480 85264
rect 439520 84872 440000 84992
rect 0 83512 480 83632
rect 439520 83512 440000 83632
rect 439520 82152 440000 82272
rect 0 81880 480 82000
rect 439520 80792 440000 80912
rect 0 80248 480 80368
rect 439520 79432 440000 79552
rect 0 78616 480 78736
rect 439520 78072 440000 78192
rect 0 76984 480 77104
rect 439520 76712 440000 76832
rect 0 75352 480 75472
rect 439520 75352 440000 75472
rect 439520 73992 440000 74112
rect 0 73720 480 73840
rect 439520 72632 440000 72752
rect 0 72088 480 72208
rect 439520 71272 440000 71392
rect 0 70456 480 70576
rect 439520 69912 440000 70032
rect 0 68824 480 68944
rect 439520 68552 440000 68672
rect 0 67192 480 67312
rect 439520 67192 440000 67312
rect 439520 65832 440000 65952
rect 0 65560 480 65680
rect 439520 64472 440000 64592
rect 0 63928 480 64048
rect 439520 63112 440000 63232
rect 0 62296 480 62416
rect 439520 61752 440000 61872
rect 0 60664 480 60784
rect 439520 60392 440000 60512
rect 0 59032 480 59152
rect 439520 59032 440000 59152
rect 439520 57672 440000 57792
rect 0 57400 480 57520
rect 439520 56312 440000 56432
rect 0 55768 480 55888
rect 439520 54952 440000 55072
rect 0 54136 480 54256
rect 439520 53592 440000 53712
rect 0 52504 480 52624
rect 439520 52232 440000 52352
rect 0 50872 480 50992
rect 439520 50872 440000 50992
rect 439520 49512 440000 49632
rect 0 49240 480 49360
rect 439520 48152 440000 48272
rect 0 47608 480 47728
rect 439520 46792 440000 46912
rect 0 45976 480 46096
rect 439520 45432 440000 45552
rect 0 44344 480 44464
rect 439520 44072 440000 44192
rect 0 42712 480 42832
rect 439520 42712 440000 42832
rect 439520 41352 440000 41472
rect 0 41080 480 41200
rect 439520 39992 440000 40112
rect 0 39448 480 39568
rect 439520 38632 440000 38752
rect 0 37816 480 37936
rect 439520 37272 440000 37392
rect 0 36184 480 36304
rect 439520 35912 440000 36032
rect 0 34552 480 34672
rect 439520 34552 440000 34672
rect 439520 33192 440000 33312
rect 0 32920 480 33040
rect 439520 31832 440000 31952
rect 0 31288 480 31408
rect 439520 30472 440000 30592
rect 0 29656 480 29776
rect 439520 29112 440000 29232
rect 0 28024 480 28144
rect 439520 27752 440000 27872
rect 0 26392 480 26512
rect 439520 26392 440000 26512
rect 439520 25032 440000 25152
rect 0 24760 480 24880
rect 439520 23672 440000 23792
rect 0 23128 480 23248
rect 439520 22312 440000 22432
rect 0 21496 480 21616
rect 439520 20952 440000 21072
rect 0 19864 480 19984
rect 439520 19592 440000 19712
rect 0 18232 480 18352
rect 439520 18232 440000 18352
rect 0 16600 480 16720
rect 0 14968 480 15088
rect 0 13336 480 13456
rect 0 11704 480 11824
rect 0 10072 480 10192
rect 0 8440 480 8560
rect 0 6808 480 6928
rect 0 5176 480 5296
rect 0 3544 480 3664
rect 0 1912 480 2032
<< obsm3 >>
rect 13 276288 439520 277541
rect 560 276008 439520 276288
rect 13 274656 439520 276008
rect 560 274376 439520 274656
rect 13 273024 439520 274376
rect 560 272744 439520 273024
rect 13 271392 439520 272744
rect 560 271112 439520 271392
rect 13 269760 439520 271112
rect 560 269480 439520 269760
rect 13 268128 439520 269480
rect 560 267848 439520 268128
rect 13 266496 439520 267848
rect 560 266216 439520 266496
rect 13 264864 439520 266216
rect 560 264584 439520 264864
rect 13 263232 439520 264584
rect 560 262952 439520 263232
rect 13 261872 439520 262952
rect 13 261600 439440 261872
rect 560 261592 439440 261600
rect 560 261320 439520 261592
rect 13 260512 439520 261320
rect 13 260232 439440 260512
rect 13 259968 439520 260232
rect 560 259688 439520 259968
rect 13 259152 439520 259688
rect 13 258872 439440 259152
rect 13 258336 439520 258872
rect 560 258056 439520 258336
rect 13 257792 439520 258056
rect 13 257512 439440 257792
rect 13 256704 439520 257512
rect 560 256432 439520 256704
rect 560 256424 439440 256432
rect 13 256152 439440 256424
rect 13 255072 439520 256152
rect 560 254792 439440 255072
rect 13 253712 439520 254792
rect 13 253440 439440 253712
rect 560 253432 439440 253440
rect 560 253160 439520 253432
rect 13 252352 439520 253160
rect 13 252072 439440 252352
rect 13 251808 439520 252072
rect 560 251528 439520 251808
rect 13 250992 439520 251528
rect 13 250712 439440 250992
rect 13 250176 439520 250712
rect 560 249896 439520 250176
rect 13 249632 439520 249896
rect 13 249352 439440 249632
rect 13 248544 439520 249352
rect 560 248272 439520 248544
rect 560 248264 439440 248272
rect 13 247992 439440 248264
rect 13 246912 439520 247992
rect 560 246632 439440 246912
rect 13 245552 439520 246632
rect 13 245280 439440 245552
rect 560 245272 439440 245280
rect 560 245000 439520 245272
rect 13 244192 439520 245000
rect 13 243912 439440 244192
rect 13 243648 439520 243912
rect 560 243368 439520 243648
rect 13 242832 439520 243368
rect 13 242552 439440 242832
rect 13 242016 439520 242552
rect 560 241736 439520 242016
rect 13 241472 439520 241736
rect 13 241192 439440 241472
rect 13 240384 439520 241192
rect 560 240112 439520 240384
rect 560 240104 439440 240112
rect 13 239832 439440 240104
rect 13 238752 439520 239832
rect 560 238472 439440 238752
rect 13 237392 439520 238472
rect 13 237120 439440 237392
rect 560 237112 439440 237120
rect 560 236840 439520 237112
rect 13 236032 439520 236840
rect 13 235752 439440 236032
rect 13 235488 439520 235752
rect 560 235208 439520 235488
rect 13 234672 439520 235208
rect 13 234392 439440 234672
rect 13 233856 439520 234392
rect 560 233576 439520 233856
rect 13 233312 439520 233576
rect 13 233032 439440 233312
rect 13 232224 439520 233032
rect 560 231952 439520 232224
rect 560 231944 439440 231952
rect 13 231672 439440 231944
rect 13 230592 439520 231672
rect 560 230312 439440 230592
rect 13 229232 439520 230312
rect 13 228960 439440 229232
rect 560 228952 439440 228960
rect 560 228680 439520 228952
rect 13 227872 439520 228680
rect 13 227592 439440 227872
rect 13 227328 439520 227592
rect 560 227048 439520 227328
rect 13 226512 439520 227048
rect 13 226232 439440 226512
rect 13 225696 439520 226232
rect 560 225416 439520 225696
rect 13 225152 439520 225416
rect 13 224872 439440 225152
rect 13 224064 439520 224872
rect 560 223792 439520 224064
rect 560 223784 439440 223792
rect 13 223512 439440 223784
rect 13 222432 439520 223512
rect 560 222152 439440 222432
rect 13 221072 439520 222152
rect 13 220800 439440 221072
rect 560 220792 439440 220800
rect 560 220520 439520 220792
rect 13 219712 439520 220520
rect 13 219432 439440 219712
rect 13 219168 439520 219432
rect 560 218888 439520 219168
rect 13 218352 439520 218888
rect 13 218072 439440 218352
rect 13 217536 439520 218072
rect 560 217256 439520 217536
rect 13 216992 439520 217256
rect 13 216712 439440 216992
rect 13 215904 439520 216712
rect 560 215632 439520 215904
rect 560 215624 439440 215632
rect 13 215352 439440 215624
rect 13 214272 439520 215352
rect 560 213992 439440 214272
rect 13 212912 439520 213992
rect 13 212640 439440 212912
rect 560 212632 439440 212640
rect 560 212360 439520 212632
rect 13 211552 439520 212360
rect 13 211272 439440 211552
rect 13 211008 439520 211272
rect 560 210728 439520 211008
rect 13 210192 439520 210728
rect 13 209912 439440 210192
rect 13 209376 439520 209912
rect 560 209096 439520 209376
rect 13 208832 439520 209096
rect 13 208552 439440 208832
rect 13 207744 439520 208552
rect 560 207472 439520 207744
rect 560 207464 439440 207472
rect 13 207192 439440 207464
rect 13 206112 439520 207192
rect 560 205832 439440 206112
rect 13 204752 439520 205832
rect 13 204480 439440 204752
rect 560 204472 439440 204480
rect 560 204200 439520 204472
rect 13 203392 439520 204200
rect 13 203112 439440 203392
rect 13 202848 439520 203112
rect 560 202568 439520 202848
rect 13 202032 439520 202568
rect 13 201752 439440 202032
rect 13 201216 439520 201752
rect 560 200936 439520 201216
rect 13 200672 439520 200936
rect 13 200392 439440 200672
rect 13 199584 439520 200392
rect 560 199312 439520 199584
rect 560 199304 439440 199312
rect 13 199032 439440 199304
rect 13 197952 439520 199032
rect 560 197672 439440 197952
rect 13 196592 439520 197672
rect 13 196320 439440 196592
rect 560 196312 439440 196320
rect 560 196040 439520 196312
rect 13 195232 439520 196040
rect 13 194952 439440 195232
rect 13 194688 439520 194952
rect 560 194408 439520 194688
rect 13 193872 439520 194408
rect 13 193592 439440 193872
rect 13 193056 439520 193592
rect 560 192776 439520 193056
rect 13 192512 439520 192776
rect 13 192232 439440 192512
rect 13 191424 439520 192232
rect 560 191152 439520 191424
rect 560 191144 439440 191152
rect 13 190872 439440 191144
rect 13 189792 439520 190872
rect 560 189512 439440 189792
rect 13 188432 439520 189512
rect 13 188160 439440 188432
rect 560 188152 439440 188160
rect 560 187880 439520 188152
rect 13 187072 439520 187880
rect 13 186792 439440 187072
rect 13 186528 439520 186792
rect 560 186248 439520 186528
rect 13 185712 439520 186248
rect 13 185432 439440 185712
rect 13 184896 439520 185432
rect 560 184616 439520 184896
rect 13 184352 439520 184616
rect 13 184072 439440 184352
rect 13 183264 439520 184072
rect 560 182992 439520 183264
rect 560 182984 439440 182992
rect 13 182712 439440 182984
rect 13 181632 439520 182712
rect 560 181352 439440 181632
rect 13 180272 439520 181352
rect 13 180000 439440 180272
rect 560 179992 439440 180000
rect 560 179720 439520 179992
rect 13 178912 439520 179720
rect 13 178632 439440 178912
rect 13 178368 439520 178632
rect 560 178088 439520 178368
rect 13 177552 439520 178088
rect 13 177272 439440 177552
rect 13 176736 439520 177272
rect 560 176456 439520 176736
rect 13 176192 439520 176456
rect 13 175912 439440 176192
rect 13 175104 439520 175912
rect 560 174832 439520 175104
rect 560 174824 439440 174832
rect 13 174552 439440 174824
rect 13 173472 439520 174552
rect 560 173192 439440 173472
rect 13 172112 439520 173192
rect 13 171840 439440 172112
rect 560 171832 439440 171840
rect 560 171560 439520 171832
rect 13 170752 439520 171560
rect 13 170472 439440 170752
rect 13 170208 439520 170472
rect 560 169928 439520 170208
rect 13 169392 439520 169928
rect 13 169112 439440 169392
rect 13 168576 439520 169112
rect 560 168296 439520 168576
rect 13 168032 439520 168296
rect 13 167752 439440 168032
rect 13 166944 439520 167752
rect 560 166672 439520 166944
rect 560 166664 439440 166672
rect 13 166392 439440 166664
rect 13 165312 439520 166392
rect 560 165032 439440 165312
rect 13 163952 439520 165032
rect 13 163680 439440 163952
rect 560 163672 439440 163680
rect 560 163400 439520 163672
rect 13 162592 439520 163400
rect 13 162312 439440 162592
rect 13 162048 439520 162312
rect 560 161768 439520 162048
rect 13 161232 439520 161768
rect 13 160952 439440 161232
rect 13 160416 439520 160952
rect 560 160136 439520 160416
rect 13 159872 439520 160136
rect 13 159592 439440 159872
rect 13 158784 439520 159592
rect 560 158512 439520 158784
rect 560 158504 439440 158512
rect 13 158232 439440 158504
rect 13 157152 439520 158232
rect 560 156872 439440 157152
rect 13 155792 439520 156872
rect 13 155520 439440 155792
rect 560 155512 439440 155520
rect 560 155240 439520 155512
rect 13 154432 439520 155240
rect 13 154152 439440 154432
rect 13 153888 439520 154152
rect 560 153608 439520 153888
rect 13 153072 439520 153608
rect 13 152792 439440 153072
rect 13 152256 439520 152792
rect 560 151976 439520 152256
rect 13 151712 439520 151976
rect 13 151432 439440 151712
rect 13 150624 439520 151432
rect 560 150352 439520 150624
rect 560 150344 439440 150352
rect 13 150072 439440 150344
rect 13 148992 439520 150072
rect 560 148712 439440 148992
rect 13 147632 439520 148712
rect 13 147360 439440 147632
rect 560 147352 439440 147360
rect 560 147080 439520 147352
rect 13 146272 439520 147080
rect 13 145992 439440 146272
rect 13 145728 439520 145992
rect 560 145448 439520 145728
rect 13 144912 439520 145448
rect 13 144632 439440 144912
rect 13 144096 439520 144632
rect 560 143816 439520 144096
rect 13 143552 439520 143816
rect 13 143272 439440 143552
rect 13 142464 439520 143272
rect 560 142192 439520 142464
rect 560 142184 439440 142192
rect 13 141912 439440 142184
rect 13 140832 439520 141912
rect 560 140552 439440 140832
rect 13 139472 439520 140552
rect 13 139200 439440 139472
rect 560 139192 439440 139200
rect 560 138920 439520 139192
rect 13 138112 439520 138920
rect 13 137832 439440 138112
rect 13 137568 439520 137832
rect 560 137288 439520 137568
rect 13 136752 439520 137288
rect 13 136472 439440 136752
rect 13 135936 439520 136472
rect 560 135656 439520 135936
rect 13 135392 439520 135656
rect 13 135112 439440 135392
rect 13 134304 439520 135112
rect 560 134032 439520 134304
rect 560 134024 439440 134032
rect 13 133752 439440 134024
rect 13 132672 439520 133752
rect 560 132392 439440 132672
rect 13 131312 439520 132392
rect 13 131040 439440 131312
rect 560 131032 439440 131040
rect 560 130760 439520 131032
rect 13 129952 439520 130760
rect 13 129672 439440 129952
rect 13 129408 439520 129672
rect 560 129128 439520 129408
rect 13 128592 439520 129128
rect 13 128312 439440 128592
rect 13 127776 439520 128312
rect 560 127496 439520 127776
rect 13 127232 439520 127496
rect 13 126952 439440 127232
rect 13 126144 439520 126952
rect 560 125872 439520 126144
rect 560 125864 439440 125872
rect 13 125592 439440 125864
rect 13 124512 439520 125592
rect 560 124232 439440 124512
rect 13 123152 439520 124232
rect 13 122880 439440 123152
rect 560 122872 439440 122880
rect 560 122600 439520 122872
rect 13 121792 439520 122600
rect 13 121512 439440 121792
rect 13 121248 439520 121512
rect 560 120968 439520 121248
rect 13 120432 439520 120968
rect 13 120152 439440 120432
rect 13 119616 439520 120152
rect 560 119336 439520 119616
rect 13 119072 439520 119336
rect 13 118792 439440 119072
rect 13 117984 439520 118792
rect 560 117712 439520 117984
rect 560 117704 439440 117712
rect 13 117432 439440 117704
rect 13 116352 439520 117432
rect 560 116072 439440 116352
rect 13 114992 439520 116072
rect 13 114720 439440 114992
rect 560 114712 439440 114720
rect 560 114440 439520 114712
rect 13 113632 439520 114440
rect 13 113352 439440 113632
rect 13 113088 439520 113352
rect 560 112808 439520 113088
rect 13 112272 439520 112808
rect 13 111992 439440 112272
rect 13 111456 439520 111992
rect 560 111176 439520 111456
rect 13 110912 439520 111176
rect 13 110632 439440 110912
rect 13 109824 439520 110632
rect 560 109552 439520 109824
rect 560 109544 439440 109552
rect 13 109272 439440 109544
rect 13 108192 439520 109272
rect 560 107912 439440 108192
rect 13 106832 439520 107912
rect 13 106560 439440 106832
rect 560 106552 439440 106560
rect 560 106280 439520 106552
rect 13 105472 439520 106280
rect 13 105192 439440 105472
rect 13 104928 439520 105192
rect 560 104648 439520 104928
rect 13 104112 439520 104648
rect 13 103832 439440 104112
rect 13 103296 439520 103832
rect 560 103016 439520 103296
rect 13 102752 439520 103016
rect 13 102472 439440 102752
rect 13 101664 439520 102472
rect 560 101392 439520 101664
rect 560 101384 439440 101392
rect 13 101112 439440 101384
rect 13 100032 439520 101112
rect 560 99752 439440 100032
rect 13 98672 439520 99752
rect 13 98400 439440 98672
rect 560 98392 439440 98400
rect 560 98120 439520 98392
rect 13 97312 439520 98120
rect 13 97032 439440 97312
rect 13 96768 439520 97032
rect 560 96488 439520 96768
rect 13 95952 439520 96488
rect 13 95672 439440 95952
rect 13 95136 439520 95672
rect 560 94856 439520 95136
rect 13 94592 439520 94856
rect 13 94312 439440 94592
rect 13 93504 439520 94312
rect 560 93232 439520 93504
rect 560 93224 439440 93232
rect 13 92952 439440 93224
rect 13 91872 439520 92952
rect 560 91592 439440 91872
rect 13 90512 439520 91592
rect 13 90240 439440 90512
rect 560 90232 439440 90240
rect 560 89960 439520 90232
rect 13 89152 439520 89960
rect 13 88872 439440 89152
rect 13 88608 439520 88872
rect 560 88328 439520 88608
rect 13 87792 439520 88328
rect 13 87512 439440 87792
rect 13 86976 439520 87512
rect 560 86696 439520 86976
rect 13 86432 439520 86696
rect 13 86152 439440 86432
rect 13 85344 439520 86152
rect 560 85072 439520 85344
rect 560 85064 439440 85072
rect 13 84792 439440 85064
rect 13 83712 439520 84792
rect 560 83432 439440 83712
rect 13 82352 439520 83432
rect 13 82080 439440 82352
rect 560 82072 439440 82080
rect 560 81800 439520 82072
rect 13 80992 439520 81800
rect 13 80712 439440 80992
rect 13 80448 439520 80712
rect 560 80168 439520 80448
rect 13 79632 439520 80168
rect 13 79352 439440 79632
rect 13 78816 439520 79352
rect 560 78536 439520 78816
rect 13 78272 439520 78536
rect 13 77992 439440 78272
rect 13 77184 439520 77992
rect 560 76912 439520 77184
rect 560 76904 439440 76912
rect 13 76632 439440 76904
rect 13 75552 439520 76632
rect 560 75272 439440 75552
rect 13 74192 439520 75272
rect 13 73920 439440 74192
rect 560 73912 439440 73920
rect 560 73640 439520 73912
rect 13 72832 439520 73640
rect 13 72552 439440 72832
rect 13 72288 439520 72552
rect 560 72008 439520 72288
rect 13 71472 439520 72008
rect 13 71192 439440 71472
rect 13 70656 439520 71192
rect 560 70376 439520 70656
rect 13 70112 439520 70376
rect 13 69832 439440 70112
rect 13 69024 439520 69832
rect 560 68752 439520 69024
rect 560 68744 439440 68752
rect 13 68472 439440 68744
rect 13 67392 439520 68472
rect 560 67112 439440 67392
rect 13 66032 439520 67112
rect 13 65760 439440 66032
rect 560 65752 439440 65760
rect 560 65480 439520 65752
rect 13 64672 439520 65480
rect 13 64392 439440 64672
rect 13 64128 439520 64392
rect 560 63848 439520 64128
rect 13 63312 439520 63848
rect 13 63032 439440 63312
rect 13 62496 439520 63032
rect 560 62216 439520 62496
rect 13 61952 439520 62216
rect 13 61672 439440 61952
rect 13 60864 439520 61672
rect 560 60592 439520 60864
rect 560 60584 439440 60592
rect 13 60312 439440 60584
rect 13 59232 439520 60312
rect 560 58952 439440 59232
rect 13 57872 439520 58952
rect 13 57600 439440 57872
rect 560 57592 439440 57600
rect 560 57320 439520 57592
rect 13 56512 439520 57320
rect 13 56232 439440 56512
rect 13 55968 439520 56232
rect 560 55688 439520 55968
rect 13 55152 439520 55688
rect 13 54872 439440 55152
rect 13 54336 439520 54872
rect 560 54056 439520 54336
rect 13 53792 439520 54056
rect 13 53512 439440 53792
rect 13 52704 439520 53512
rect 560 52432 439520 52704
rect 560 52424 439440 52432
rect 13 52152 439440 52424
rect 13 51072 439520 52152
rect 560 50792 439440 51072
rect 13 49712 439520 50792
rect 13 49440 439440 49712
rect 560 49432 439440 49440
rect 560 49160 439520 49432
rect 13 48352 439520 49160
rect 13 48072 439440 48352
rect 13 47808 439520 48072
rect 560 47528 439520 47808
rect 13 46992 439520 47528
rect 13 46712 439440 46992
rect 13 46176 439520 46712
rect 560 45896 439520 46176
rect 13 45632 439520 45896
rect 13 45352 439440 45632
rect 13 44544 439520 45352
rect 560 44272 439520 44544
rect 560 44264 439440 44272
rect 13 43992 439440 44264
rect 13 42912 439520 43992
rect 560 42632 439440 42912
rect 13 41552 439520 42632
rect 13 41280 439440 41552
rect 560 41272 439440 41280
rect 560 41000 439520 41272
rect 13 40192 439520 41000
rect 13 39912 439440 40192
rect 13 39648 439520 39912
rect 560 39368 439520 39648
rect 13 38832 439520 39368
rect 13 38552 439440 38832
rect 13 38016 439520 38552
rect 560 37736 439520 38016
rect 13 37472 439520 37736
rect 13 37192 439440 37472
rect 13 36384 439520 37192
rect 560 36112 439520 36384
rect 560 36104 439440 36112
rect 13 35832 439440 36104
rect 13 34752 439520 35832
rect 560 34472 439440 34752
rect 13 33392 439520 34472
rect 13 33120 439440 33392
rect 560 33112 439440 33120
rect 560 32840 439520 33112
rect 13 32032 439520 32840
rect 13 31752 439440 32032
rect 13 31488 439520 31752
rect 560 31208 439520 31488
rect 13 30672 439520 31208
rect 13 30392 439440 30672
rect 13 29856 439520 30392
rect 560 29576 439520 29856
rect 13 29312 439520 29576
rect 13 29032 439440 29312
rect 13 28224 439520 29032
rect 560 27952 439520 28224
rect 560 27944 439440 27952
rect 13 27672 439440 27944
rect 13 26592 439520 27672
rect 560 26312 439440 26592
rect 13 25232 439520 26312
rect 13 24960 439440 25232
rect 560 24952 439440 24960
rect 560 24680 439520 24952
rect 13 23872 439520 24680
rect 13 23592 439440 23872
rect 13 23328 439520 23592
rect 560 23048 439520 23328
rect 13 22512 439520 23048
rect 13 22232 439440 22512
rect 13 21696 439520 22232
rect 560 21416 439520 21696
rect 13 21152 439520 21416
rect 13 20872 439440 21152
rect 13 20064 439520 20872
rect 560 19792 439520 20064
rect 560 19784 439440 19792
rect 13 19512 439440 19784
rect 13 18432 439520 19512
rect 560 18152 439440 18432
rect 13 16800 439520 18152
rect 560 16520 439520 16800
rect 13 15168 439520 16520
rect 560 14888 439520 15168
rect 13 13536 439520 14888
rect 560 13256 439520 13536
rect 13 11904 439520 13256
rect 560 11624 439520 11904
rect 13 10272 439520 11624
rect 560 9992 439520 10272
rect 13 8640 439520 9992
rect 560 8360 439520 8640
rect 13 7008 439520 8360
rect 560 6728 439520 7008
rect 13 5376 439520 6728
rect 560 5096 439520 5376
rect 13 3744 439520 5096
rect 560 3464 439520 3744
rect 13 2143 439520 3464
<< metal4 >>
rect 1794 2128 2414 277488
rect 2814 2128 3434 277488
rect 7794 2128 8414 277488
rect 8814 2128 9434 277488
rect 13794 2128 14414 277488
rect 14814 2128 15434 277488
rect 19794 165388 20414 277488
rect 20814 165328 21434 277488
rect 25794 165388 26414 277488
rect 26814 165328 27434 277488
rect 31794 165388 32414 277488
rect 32814 165328 33434 277488
rect 37794 165388 38414 277488
rect 38814 165328 39434 277488
rect 43794 165388 44414 277488
rect 44814 165328 45434 277488
rect 49794 165388 50414 277488
rect 50814 165373 51434 277488
rect 55794 165388 56414 277488
rect 56814 165328 57434 277488
rect 61794 165388 62414 277488
rect 62814 165373 63434 277488
rect 67794 165388 68414 277488
rect 68814 165328 69434 277488
rect 73794 165388 74414 277488
rect 74814 165328 75434 277488
rect 79794 165388 80414 277488
rect 80814 165373 81434 277488
rect 85794 165388 86414 277488
rect 86814 165328 87434 277488
rect 91794 165388 92414 277488
rect 92814 165328 93434 277488
rect 97794 165388 98414 277488
rect 98814 165328 99434 277488
rect 103794 165388 104414 277488
rect 104814 165328 105434 277488
rect 109794 165388 110414 277488
rect 110814 165373 111434 277488
rect 115794 165388 116414 277488
rect 116814 165328 117434 277488
rect 121794 165388 122414 277488
rect 122814 165373 123434 277488
rect 127794 165388 128414 277488
rect 128814 165328 129434 277488
rect 133794 165388 134414 277488
rect 134814 165328 135434 277488
rect 139794 165388 140414 277488
rect 140814 165328 141434 277488
rect 145794 165388 146414 277488
rect 146814 165328 147434 277488
rect 151794 165388 152414 277488
rect 152814 165328 153434 277488
rect 157794 165388 158414 277488
rect 19794 2128 20414 77920
rect 20814 2128 21434 77920
rect 25794 2128 26414 77920
rect 26814 2128 27434 77920
rect 31794 2128 32414 77920
rect 32814 2128 33434 77920
rect 37794 2128 38414 77920
rect 38814 2128 39434 77920
rect 43794 2128 44414 77920
rect 44814 2128 45434 77920
rect 49794 2128 50414 77920
rect 50814 2128 51434 77920
rect 55794 2128 56414 77920
rect 56814 2128 57434 77920
rect 61794 2128 62414 77920
rect 62814 2128 63434 77920
rect 67794 2128 68414 77920
rect 68814 2128 69434 77920
rect 73794 2128 74414 77920
rect 74814 2128 75434 77920
rect 79794 2128 80414 77920
rect 80814 2128 81434 77920
rect 85794 2128 86414 77920
rect 86814 2128 87434 77920
rect 91794 2128 92414 77920
rect 92814 2128 93434 77920
rect 97794 2128 98414 77920
rect 98814 2128 99434 77920
rect 103794 2128 104414 77920
rect 104814 2128 105434 77920
rect 109794 2128 110414 77920
rect 110814 2128 111434 77920
rect 115794 2128 116414 77920
rect 116814 2128 117434 77920
rect 121794 2128 122414 77920
rect 122814 2128 123434 77920
rect 127794 2128 128414 77920
rect 128814 2128 129434 77920
rect 133794 2128 134414 77920
rect 134814 2128 135434 77920
rect 139794 2128 140414 77920
rect 140814 2128 141434 77920
rect 145794 2128 146414 77920
rect 146814 2128 147434 77920
rect 151794 2128 152414 77920
rect 152814 2128 153434 77920
rect 157794 2128 158414 77920
rect 158814 2128 159434 277488
rect 163794 2128 164414 277488
rect 164814 2128 165434 277488
rect 169794 2128 170414 277488
rect 170814 2128 171434 277488
rect 175794 2128 176414 277488
rect 176814 2128 177434 277488
rect 181794 2128 182414 277488
rect 182814 2128 183434 277488
rect 187794 2128 188414 277488
rect 188814 2128 189434 277488
rect 193794 2128 194414 277488
rect 194814 2128 195434 277488
rect 199794 2128 200414 277488
rect 200814 2128 201434 277488
rect 205794 69040 206414 277488
rect 206814 69080 207434 277488
rect 211794 69040 212414 277488
rect 212814 69080 213434 277488
rect 217794 69040 218414 277488
rect 218814 69080 219434 277488
rect 223794 69040 224414 277488
rect 224814 69080 225434 277488
rect 205794 2128 206414 49920
rect 206814 2128 207434 49920
rect 211794 2128 212414 49920
rect 212814 2128 213434 49920
rect 217794 2128 218414 49920
rect 218814 2128 219434 49920
rect 223794 2128 224414 49920
rect 224814 2128 225434 49920
rect 229794 2128 230414 277488
rect 230814 2128 231434 277488
rect 235794 2128 236414 277488
rect 236814 2128 237434 277488
rect 241794 2128 242414 277488
rect 242814 2128 243434 277488
rect 247794 2128 248414 277488
rect 248814 2128 249434 277488
rect 253794 2128 254414 277488
rect 254814 2128 255434 277488
rect 259794 2128 260414 277488
rect 260814 2128 261434 277488
rect 265794 2128 266414 277488
rect 266814 2128 267434 277488
rect 271794 2128 272414 277488
rect 272814 2128 273434 277488
rect 277794 165388 278414 277488
rect 278814 165328 279434 277488
rect 283794 165388 284414 277488
rect 284814 165328 285434 277488
rect 289794 165388 290414 277488
rect 290814 165328 291434 277488
rect 295794 165388 296414 277488
rect 296814 165328 297434 277488
rect 301794 165388 302414 277488
rect 302814 165328 303434 277488
rect 307794 165388 308414 277488
rect 308814 165328 309434 277488
rect 313794 165388 314414 277488
rect 314814 165328 315434 277488
rect 319794 165388 320414 277488
rect 320814 165373 321434 277488
rect 325794 165388 326414 277488
rect 326814 165328 327434 277488
rect 331794 165388 332414 277488
rect 332814 165328 333434 277488
rect 337794 165388 338414 277488
rect 338814 165328 339434 277488
rect 343794 165388 344414 277488
rect 344814 165328 345434 277488
rect 349794 165388 350414 277488
rect 350814 165373 351434 277488
rect 355794 165388 356414 277488
rect 356814 165328 357434 277488
rect 361794 165388 362414 277488
rect 362814 165373 363434 277488
rect 367794 165388 368414 277488
rect 368814 165328 369434 277488
rect 373794 165388 374414 277488
rect 374814 165328 375434 277488
rect 379794 165388 380414 277488
rect 380814 165373 381434 277488
rect 385794 165388 386414 277488
rect 386814 165328 387434 277488
rect 391794 165388 392414 277488
rect 392814 165328 393434 277488
rect 397794 165388 398414 277488
rect 398814 165328 399434 277488
rect 403794 165388 404414 277488
rect 404814 165328 405434 277488
rect 409794 165388 410414 277488
rect 410814 165373 411434 277488
rect 415794 165388 416414 277488
rect 416814 165328 417434 277488
rect 277794 2128 278414 77920
rect 278814 2128 279434 77920
rect 283794 2128 284414 77920
rect 284814 2128 285434 77920
rect 289794 2128 290414 77920
rect 290814 2128 291434 77920
rect 295794 2128 296414 77920
rect 296814 2128 297434 77920
rect 301794 2128 302414 77920
rect 302814 2128 303434 77920
rect 307794 2128 308414 77920
rect 308814 2128 309434 77920
rect 313794 2128 314414 77920
rect 314814 2128 315434 77920
rect 319794 2128 320414 77920
rect 320814 2128 321434 77920
rect 325794 2128 326414 77920
rect 326814 2128 327434 77920
rect 331794 2128 332414 77920
rect 332814 2128 333434 77920
rect 337794 2128 338414 77920
rect 338814 2128 339434 77920
rect 343794 2128 344414 77920
rect 344814 2128 345434 77920
rect 349794 2128 350414 77920
rect 350814 2128 351434 77920
rect 355794 2128 356414 77920
rect 356814 2128 357434 77920
rect 361794 2128 362414 77920
rect 362814 2128 363434 77920
rect 367794 2128 368414 77920
rect 368814 2128 369434 77920
rect 373794 2128 374414 77920
rect 374814 2128 375434 77920
rect 379794 2128 380414 77920
rect 380814 2128 381434 77920
rect 385794 2128 386414 77920
rect 386814 2128 387434 77920
rect 391794 2128 392414 77920
rect 392814 2128 393434 77920
rect 397794 2128 398414 77920
rect 398814 2128 399434 77920
rect 403794 2128 404414 77920
rect 404814 2128 405434 77920
rect 409794 2128 410414 77920
rect 410814 2128 411434 77920
rect 415794 2128 416414 77920
rect 416814 2128 417434 77920
rect 421794 2128 422414 277488
rect 422814 2128 423434 277488
rect 427794 2128 428414 277488
rect 428814 2128 429434 277488
rect 433794 2128 434414 277488
rect 434814 2128 435434 277488
<< obsm4 >>
rect 4291 13771 7714 270605
rect 8494 13771 8734 270605
rect 9514 13771 13714 270605
rect 14494 13771 14734 270605
rect 15514 165308 19714 270605
rect 20494 165308 20734 270605
rect 15514 165248 20734 165308
rect 21514 165308 25714 270605
rect 26494 165308 26734 270605
rect 21514 165248 26734 165308
rect 27514 165308 31714 270605
rect 32494 165308 32734 270605
rect 27514 165248 32734 165308
rect 33514 165308 37714 270605
rect 38494 165308 38734 270605
rect 33514 165248 38734 165308
rect 39514 165308 43714 270605
rect 44494 165308 44734 270605
rect 39514 165248 44734 165308
rect 45514 165308 49714 270605
rect 50494 165308 50734 270605
rect 45514 165293 50734 165308
rect 51514 165308 55714 270605
rect 56494 165308 56734 270605
rect 51514 165293 56734 165308
rect 45514 165248 56734 165293
rect 57514 165308 61714 270605
rect 62494 165308 62734 270605
rect 57514 165293 62734 165308
rect 63514 165308 67714 270605
rect 68494 165308 68734 270605
rect 63514 165293 68734 165308
rect 57514 165248 68734 165293
rect 69514 165308 73714 270605
rect 74494 165308 74734 270605
rect 69514 165248 74734 165308
rect 75514 165308 79714 270605
rect 80494 165308 80734 270605
rect 75514 165293 80734 165308
rect 81514 165308 85714 270605
rect 86494 165308 86734 270605
rect 81514 165293 86734 165308
rect 75514 165248 86734 165293
rect 87514 165308 91714 270605
rect 92494 165308 92734 270605
rect 87514 165248 92734 165308
rect 93514 165308 97714 270605
rect 98494 165308 98734 270605
rect 93514 165248 98734 165308
rect 99514 165308 103714 270605
rect 104494 165308 104734 270605
rect 99514 165248 104734 165308
rect 105514 165308 109714 270605
rect 110494 165308 110734 270605
rect 105514 165293 110734 165308
rect 111514 165308 115714 270605
rect 116494 165308 116734 270605
rect 111514 165293 116734 165308
rect 105514 165248 116734 165293
rect 117514 165308 121714 270605
rect 122494 165308 122734 270605
rect 117514 165293 122734 165308
rect 123514 165308 127714 270605
rect 128494 165308 128734 270605
rect 123514 165293 128734 165308
rect 117514 165248 128734 165293
rect 129514 165308 133714 270605
rect 134494 165308 134734 270605
rect 129514 165248 134734 165308
rect 135514 165308 139714 270605
rect 140494 165308 140734 270605
rect 135514 165248 140734 165308
rect 141514 165308 145714 270605
rect 146494 165308 146734 270605
rect 141514 165248 146734 165308
rect 147514 165308 151714 270605
rect 152494 165308 152734 270605
rect 147514 165248 152734 165308
rect 153514 165308 157714 270605
rect 158494 165308 158734 270605
rect 153514 165248 158734 165308
rect 15514 78000 158734 165248
rect 15514 13771 19714 78000
rect 20494 13771 20734 78000
rect 21514 13771 25714 78000
rect 26494 13771 26734 78000
rect 27514 13771 31714 78000
rect 32494 13771 32734 78000
rect 33514 13771 37714 78000
rect 38494 13771 38734 78000
rect 39514 13771 43714 78000
rect 44494 13771 44734 78000
rect 45514 13771 49714 78000
rect 50494 13771 50734 78000
rect 51514 13771 55714 78000
rect 56494 13771 56734 78000
rect 57514 13771 61714 78000
rect 62494 13771 62734 78000
rect 63514 13771 67714 78000
rect 68494 13771 68734 78000
rect 69514 13771 73714 78000
rect 74494 13771 74734 78000
rect 75514 13771 79714 78000
rect 80494 13771 80734 78000
rect 81514 13771 85714 78000
rect 86494 13771 86734 78000
rect 87514 13771 91714 78000
rect 92494 13771 92734 78000
rect 93514 13771 97714 78000
rect 98494 13771 98734 78000
rect 99514 13771 103714 78000
rect 104494 13771 104734 78000
rect 105514 13771 109714 78000
rect 110494 13771 110734 78000
rect 111514 13771 115714 78000
rect 116494 13771 116734 78000
rect 117514 13771 121714 78000
rect 122494 13771 122734 78000
rect 123514 13771 127714 78000
rect 128494 13771 128734 78000
rect 129514 13771 133714 78000
rect 134494 13771 134734 78000
rect 135514 13771 139714 78000
rect 140494 13771 140734 78000
rect 141514 13771 145714 78000
rect 146494 13771 146734 78000
rect 147514 13771 151714 78000
rect 152494 13771 152734 78000
rect 153514 13771 157714 78000
rect 158494 13771 158734 78000
rect 159514 13771 163714 270605
rect 164494 13771 164734 270605
rect 165514 13771 169714 270605
rect 170494 13771 170734 270605
rect 171514 13771 175714 270605
rect 176494 13771 176734 270605
rect 177514 13771 181714 270605
rect 182494 13771 182734 270605
rect 183514 13771 187714 270605
rect 188494 13771 188734 270605
rect 189514 13771 193714 270605
rect 194494 13771 194734 270605
rect 195514 13771 199714 270605
rect 200494 13771 200734 270605
rect 201514 68960 205714 270605
rect 206494 69000 206734 270605
rect 207514 69000 211714 270605
rect 206494 68960 211714 69000
rect 212494 69000 212734 270605
rect 213514 69000 217714 270605
rect 212494 68960 217714 69000
rect 218494 69000 218734 270605
rect 219514 69000 223714 270605
rect 218494 68960 223714 69000
rect 224494 69000 224734 270605
rect 225514 69000 229714 270605
rect 224494 68960 229714 69000
rect 201514 50000 229714 68960
rect 201514 13771 205714 50000
rect 206494 13771 206734 50000
rect 207514 13771 211714 50000
rect 212494 13771 212734 50000
rect 213514 13771 217714 50000
rect 218494 13771 218734 50000
rect 219514 13771 223714 50000
rect 224494 13771 224734 50000
rect 225514 13771 229714 50000
rect 230494 13771 230734 270605
rect 231514 13771 235714 270605
rect 236494 13771 236734 270605
rect 237514 13771 241714 270605
rect 242494 13771 242734 270605
rect 243514 13771 247714 270605
rect 248494 13771 248734 270605
rect 249514 13771 253714 270605
rect 254494 13771 254734 270605
rect 255514 13771 259714 270605
rect 260494 13771 260734 270605
rect 261514 13771 265714 270605
rect 266494 13771 266734 270605
rect 267514 13771 271714 270605
rect 272494 13771 272734 270605
rect 273514 165308 277714 270605
rect 278494 165308 278734 270605
rect 273514 165248 278734 165308
rect 279514 165308 283714 270605
rect 284494 165308 284734 270605
rect 279514 165248 284734 165308
rect 285514 165308 289714 270605
rect 290494 165308 290734 270605
rect 285514 165248 290734 165308
rect 291514 165308 295714 270605
rect 296494 165308 296734 270605
rect 291514 165248 296734 165308
rect 297514 165308 301714 270605
rect 302494 165308 302734 270605
rect 297514 165248 302734 165308
rect 303514 165308 307714 270605
rect 308494 165308 308734 270605
rect 303514 165248 308734 165308
rect 309514 165308 313714 270605
rect 314494 165308 314734 270605
rect 309514 165248 314734 165308
rect 315514 165308 319714 270605
rect 320494 165308 320734 270605
rect 315514 165293 320734 165308
rect 321514 165308 325714 270605
rect 326494 165308 326734 270605
rect 321514 165293 326734 165308
rect 315514 165248 326734 165293
rect 327514 165308 331714 270605
rect 332494 165308 332734 270605
rect 327514 165248 332734 165308
rect 333514 165308 337714 270605
rect 338494 165308 338734 270605
rect 333514 165248 338734 165308
rect 339514 165308 343714 270605
rect 344494 165308 344734 270605
rect 339514 165248 344734 165308
rect 345514 165308 349714 270605
rect 350494 165308 350734 270605
rect 345514 165293 350734 165308
rect 351514 165308 355714 270605
rect 356494 165308 356734 270605
rect 351514 165293 356734 165308
rect 345514 165248 356734 165293
rect 357514 165308 361714 270605
rect 362494 165308 362734 270605
rect 357514 165293 362734 165308
rect 363514 165308 367714 270605
rect 368494 165308 368734 270605
rect 363514 165293 368734 165308
rect 357514 165248 368734 165293
rect 369514 165308 373714 270605
rect 374494 165308 374734 270605
rect 369514 165248 374734 165308
rect 375514 165308 379714 270605
rect 380494 165308 380734 270605
rect 375514 165293 380734 165308
rect 381514 165308 385714 270605
rect 386494 165308 386734 270605
rect 381514 165293 386734 165308
rect 375514 165248 386734 165293
rect 387514 165308 391714 270605
rect 392494 165308 392734 270605
rect 387514 165248 392734 165308
rect 393514 165308 397714 270605
rect 398494 165308 398734 270605
rect 393514 165248 398734 165308
rect 399514 165308 403714 270605
rect 404494 165308 404734 270605
rect 399514 165248 404734 165308
rect 405514 165308 409714 270605
rect 410494 165308 410734 270605
rect 405514 165293 410734 165308
rect 411514 165308 415714 270605
rect 416494 165308 416734 270605
rect 411514 165293 416734 165308
rect 405514 165248 416734 165293
rect 417514 165248 421714 270605
rect 273514 78000 421714 165248
rect 273514 13771 277714 78000
rect 278494 13771 278734 78000
rect 279514 13771 283714 78000
rect 284494 13771 284734 78000
rect 285514 13771 289714 78000
rect 290494 13771 290734 78000
rect 291514 13771 295714 78000
rect 296494 13771 296734 78000
rect 297514 13771 301714 78000
rect 302494 13771 302734 78000
rect 303514 13771 307714 78000
rect 308494 13771 308734 78000
rect 309514 13771 313714 78000
rect 314494 13771 314734 78000
rect 315514 13771 319714 78000
rect 320494 13771 320734 78000
rect 321514 13771 325714 78000
rect 326494 13771 326734 78000
rect 327514 13771 331714 78000
rect 332494 13771 332734 78000
rect 333514 13771 337714 78000
rect 338494 13771 338734 78000
rect 339514 13771 343714 78000
rect 344494 13771 344734 78000
rect 345514 13771 349714 78000
rect 350494 13771 350734 78000
rect 351514 13771 355714 78000
rect 356494 13771 356734 78000
rect 357514 13771 361714 78000
rect 362494 13771 362734 78000
rect 363514 13771 367714 78000
rect 368494 13771 368734 78000
rect 369514 13771 373714 78000
rect 374494 13771 374734 78000
rect 375514 13771 379714 78000
rect 380494 13771 380734 78000
rect 381514 13771 385714 78000
rect 386494 13771 386734 78000
rect 387514 13771 391714 78000
rect 392494 13771 392734 78000
rect 393514 13771 397714 78000
rect 398494 13771 398734 78000
rect 399514 13771 403714 78000
rect 404494 13771 404734 78000
rect 405514 13771 409714 78000
rect 410494 13771 410734 78000
rect 411514 13771 415714 78000
rect 416494 13771 416734 78000
rect 417514 13771 421714 78000
rect 422494 13771 422734 270605
rect 423514 13771 427714 270605
rect 428494 13771 428734 270605
rect 429514 13771 433714 270605
rect 434494 13771 434734 270605
rect 435514 13771 436757 270605
<< metal5 >>
rect 1056 275886 438888 276506
rect 1056 274866 438888 275486
rect 1056 267886 438888 268506
rect 1056 266866 438888 267486
rect 1056 259886 438888 260506
rect 1056 258866 438888 259486
rect 1056 251886 438888 252506
rect 1056 250866 438888 251486
rect 1056 243886 438888 244506
rect 1056 242866 438888 243486
rect 1056 235886 438888 236506
rect 1056 234866 438888 235486
rect 1056 227886 438888 228506
rect 1056 226866 438888 227486
rect 1056 219886 438888 220506
rect 1056 218866 438888 219486
rect 1056 211886 438888 212506
rect 1056 210866 438888 211486
rect 1056 203886 438888 204506
rect 1056 202866 438888 203486
rect 1056 195886 438888 196506
rect 1056 194866 438888 195486
rect 1056 187886 438888 188506
rect 1056 186866 438888 187486
rect 1056 179886 438888 180506
rect 1056 178866 438888 179486
rect 1056 171886 438888 172506
rect 1056 170866 438888 171486
rect 1056 163886 438888 164506
rect 1056 162866 438888 163486
rect 1056 155886 438888 156506
rect 1056 154866 438888 155486
rect 1056 147886 438888 148506
rect 1056 146866 438888 147486
rect 1056 139886 438888 140506
rect 1056 138866 438888 139486
rect 1056 131886 438888 132506
rect 1056 130866 438888 131486
rect 1056 123886 438888 124506
rect 1056 122866 438888 123486
rect 1056 115886 438888 116506
rect 1056 114866 438888 115486
rect 1056 107886 438888 108506
rect 1056 106866 438888 107486
rect 1056 99886 438888 100506
rect 1056 98866 438888 99486
rect 1056 91886 438888 92506
rect 1056 90866 438888 91486
rect 1056 83886 438888 84506
rect 1056 82866 438888 83486
rect 1056 75886 438888 76506
rect 1056 74866 438888 75486
rect 1056 67886 438888 68506
rect 1056 66866 438888 67486
rect 1056 59886 438888 60506
rect 1056 58866 438888 59486
rect 1056 51886 438888 52506
rect 1056 50866 438888 51486
rect 1056 43886 438888 44506
rect 1056 42866 438888 43486
rect 1056 35886 438888 36506
rect 1056 34866 438888 35486
rect 1056 27886 438888 28506
rect 1056 26866 438888 27486
rect 1056 19886 438888 20506
rect 1056 18866 438888 19486
rect 1056 11886 438888 12506
rect 1056 10866 438888 11486
rect 1056 3886 438888 4506
rect 1056 2866 438888 3486
<< obsm5 >>
rect 10788 172826 424188 177980
rect 10788 164826 424188 170546
rect 10788 156826 424188 162546
rect 10788 148826 424188 154546
rect 10788 140826 424188 146546
rect 10788 132826 424188 138546
rect 10788 124826 424188 130546
rect 10788 116826 424188 122546
rect 10788 108826 424188 114546
rect 10788 100826 424188 106546
rect 10788 92826 424188 98546
rect 10788 84826 424188 90546
rect 10788 76826 424188 82546
rect 10788 68826 424188 74546
rect 10788 60826 424188 66546
rect 10788 55940 424188 58546
<< labels >>
rlabel metal5 s 1056 275886 438888 276506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 267886 438888 268506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 259886 438888 260506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 251886 438888 252506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 243886 438888 244506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 235886 438888 236506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 227886 438888 228506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 219886 438888 220506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 211886 438888 212506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 203886 438888 204506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 195886 438888 196506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 187886 438888 188506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 179886 438888 180506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 171886 438888 172506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 163886 438888 164506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 155886 438888 156506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 147886 438888 148506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 139886 438888 140506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 131886 438888 132506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 123886 438888 124506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 115886 438888 116506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 107886 438888 108506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 99886 438888 100506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 91886 438888 92506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 83886 438888 84506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 75886 438888 76506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 67886 438888 68506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 59886 438888 60506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 51886 438888 52506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 43886 438888 44506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 35886 438888 36506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 27886 438888 28506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 19886 438888 20506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 11886 438888 12506 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 3886 438888 4506 6 VGND
port 1 nsew ground default
rlabel metal4 s 434814 2128 435434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 428814 2128 429434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 422814 2128 423434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 416814 165328 417434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 416814 2128 417434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 410814 165373 411434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 410814 2128 411434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 404814 165328 405434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 404814 2128 405434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 398814 165328 399434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 398814 2128 399434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 392814 165328 393434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 392814 2128 393434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 386814 165328 387434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 386814 2128 387434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 380814 165373 381434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 380814 2128 381434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 374814 165328 375434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 374814 2128 375434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 368814 165328 369434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 368814 2128 369434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 362814 165373 363434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 362814 2128 363434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 356814 165328 357434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 356814 2128 357434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 350814 165373 351434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 350814 2128 351434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 344814 165328 345434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 344814 2128 345434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 338814 165328 339434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 338814 2128 339434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 332814 165328 333434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 332814 2128 333434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 326814 165328 327434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 326814 2128 327434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 320814 165373 321434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 320814 2128 321434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 314814 165328 315434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 314814 2128 315434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 308814 165328 309434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 308814 2128 309434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 302814 165328 303434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 302814 2128 303434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 296814 165328 297434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 296814 2128 297434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 290814 165328 291434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 290814 2128 291434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 284814 165328 285434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 284814 2128 285434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 278814 165328 279434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 278814 2128 279434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 272814 2128 273434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 266814 2128 267434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 260814 2128 261434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 254814 2128 255434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 248814 2128 249434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 242814 2128 243434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 236814 2128 237434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 230814 2128 231434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 224814 69080 225434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 224814 2128 225434 49920 6 VGND
port 1 nsew ground default
rlabel metal4 s 218814 69080 219434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 218814 2128 219434 49920 6 VGND
port 1 nsew ground default
rlabel metal4 s 212814 69080 213434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 212814 2128 213434 49920 6 VGND
port 1 nsew ground default
rlabel metal4 s 206814 69080 207434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 206814 2128 207434 49920 6 VGND
port 1 nsew ground default
rlabel metal4 s 200814 2128 201434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 194814 2128 195434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 188814 2128 189434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 182814 2128 183434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 176814 2128 177434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 170814 2128 171434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 164814 2128 165434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 158814 2128 159434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 152814 165328 153434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 152814 2128 153434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 146814 165328 147434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 146814 2128 147434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 140814 165328 141434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 140814 2128 141434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 134814 165328 135434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 134814 2128 135434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 128814 165328 129434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 128814 2128 129434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 122814 165373 123434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 122814 2128 123434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 116814 165328 117434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 116814 2128 117434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 110814 165373 111434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 110814 2128 111434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 104814 165328 105434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 104814 2128 105434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 98814 165328 99434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 98814 2128 99434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 92814 165328 93434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 92814 2128 93434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 86814 165328 87434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 86814 2128 87434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 80814 165373 81434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 80814 2128 81434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 74814 165328 75434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 74814 2128 75434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 68814 165328 69434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 68814 2128 69434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 62814 165373 63434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 62814 2128 63434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 56814 165328 57434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 56814 2128 57434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 50814 165373 51434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 50814 2128 51434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 44814 165328 45434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 44814 2128 45434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 38814 165328 39434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 38814 2128 39434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 32814 165328 33434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 32814 2128 33434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 26814 165328 27434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 26814 2128 27434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 20814 165328 21434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 20814 2128 21434 77920 6 VGND
port 1 nsew ground default
rlabel metal4 s 14814 2128 15434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 8814 2128 9434 277488 6 VGND
port 1 nsew ground default
rlabel metal4 s 2814 2128 3434 277488 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 274866 438888 275486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 266866 438888 267486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 258866 438888 259486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 250866 438888 251486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 242866 438888 243486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 234866 438888 235486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 226866 438888 227486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 218866 438888 219486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 210866 438888 211486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 202866 438888 203486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 194866 438888 195486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 186866 438888 187486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 178866 438888 179486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 170866 438888 171486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 162866 438888 163486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 154866 438888 155486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 146866 438888 147486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 138866 438888 139486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 130866 438888 131486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 122866 438888 123486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 114866 438888 115486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 106866 438888 107486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 98866 438888 99486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 90866 438888 91486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 82866 438888 83486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 74866 438888 75486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 66866 438888 67486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 58866 438888 59486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 50866 438888 51486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 42866 438888 43486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 34866 438888 35486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 26866 438888 27486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 18866 438888 19486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 10866 438888 11486 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 2866 438888 3486 6 VPWR
port 2 nsew power default
rlabel metal4 s 433794 2128 434414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 427794 2128 428414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 421794 2128 422414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 415794 165388 416414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 415794 2128 416414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 409794 165388 410414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 409794 2128 410414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 403794 165388 404414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 403794 2128 404414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 397794 165388 398414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 397794 2128 398414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 391794 165388 392414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 391794 2128 392414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 385794 165388 386414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 385794 2128 386414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 379794 165388 380414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 379794 2128 380414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 373794 165388 374414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 373794 2128 374414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 367794 165388 368414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 367794 2128 368414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 361794 165388 362414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 361794 2128 362414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 355794 165388 356414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 355794 2128 356414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 349794 165388 350414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 349794 2128 350414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 343794 165388 344414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 343794 2128 344414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 337794 165388 338414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 337794 2128 338414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 331794 165388 332414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 331794 2128 332414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 325794 165388 326414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 325794 2128 326414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 319794 165388 320414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 319794 2128 320414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 313794 165388 314414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 313794 2128 314414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 307794 165388 308414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 307794 2128 308414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 301794 165388 302414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 301794 2128 302414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 295794 165388 296414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 295794 2128 296414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 289794 165388 290414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 289794 2128 290414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 283794 165388 284414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 283794 2128 284414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 277794 165388 278414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 277794 2128 278414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 271794 2128 272414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 265794 2128 266414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 259794 2128 260414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 253794 2128 254414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 247794 2128 248414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 241794 2128 242414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 235794 2128 236414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 229794 2128 230414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 223794 69040 224414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 223794 2128 224414 49920 6 VPWR
port 2 nsew power default
rlabel metal4 s 217794 69040 218414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 217794 2128 218414 49920 6 VPWR
port 2 nsew power default
rlabel metal4 s 211794 69040 212414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 211794 2128 212414 49920 6 VPWR
port 2 nsew power default
rlabel metal4 s 205794 69040 206414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 205794 2128 206414 49920 6 VPWR
port 2 nsew power default
rlabel metal4 s 199794 2128 200414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 193794 2128 194414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 187794 2128 188414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 181794 2128 182414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 175794 2128 176414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 169794 2128 170414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 163794 2128 164414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 157794 165388 158414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 157794 2128 158414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 151794 165388 152414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 151794 2128 152414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 145794 165388 146414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 145794 2128 146414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 139794 165388 140414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 139794 2128 140414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 133794 165388 134414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 133794 2128 134414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 127794 165388 128414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 127794 2128 128414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 121794 165388 122414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 121794 2128 122414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 115794 165388 116414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 115794 2128 116414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 109794 165388 110414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 109794 2128 110414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 103794 165388 104414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 103794 2128 104414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 97794 165388 98414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 97794 2128 98414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 91794 165388 92414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 91794 2128 92414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 85794 165388 86414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 85794 2128 86414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 79794 165388 80414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 79794 2128 80414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 73794 165388 74414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 73794 2128 74414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 67794 165388 68414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 67794 2128 68414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 61794 165388 62414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 61794 2128 62414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 55794 165388 56414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 55794 2128 56414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 49794 165388 50414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 49794 2128 50414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 43794 165388 44414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 43794 2128 44414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 37794 165388 38414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 37794 2128 38414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 31794 165388 32414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 31794 2128 32414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 25794 165388 26414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 25794 2128 26414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 19794 165388 20414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 19794 2128 20414 77920 6 VPWR
port 2 nsew power default
rlabel metal4 s 13794 2128 14414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 7794 2128 8414 277488 6 VPWR
port 2 nsew power default
rlabel metal4 s 1794 2128 2414 277488 6 VPWR
port 2 nsew power default
rlabel metal3 s 439520 22312 440000 22432 6 gpio_dm0[0]
port 3 nsew
rlabel metal3 s 439520 185512 440000 185632 6 gpio_dm0[10]
port 4 nsew
rlabel metal3 s 439520 201832 440000 201952 6 gpio_dm0[11]
port 5 nsew
rlabel metal3 s 439520 218152 440000 218272 6 gpio_dm0[12]
port 6 nsew
rlabel metal3 s 439520 234472 440000 234592 6 gpio_dm0[13]
port 7 nsew
rlabel metal3 s 439520 250792 440000 250912 6 gpio_dm0[14]
port 8 nsew
rlabel metal2 s 424322 279520 424378 280000 6 gpio_dm0[15]
port 9 nsew
rlabel metal2 s 375746 279520 375802 280000 6 gpio_dm0[16]
port 10 nsew
rlabel metal2 s 327170 279520 327226 280000 6 gpio_dm0[17]
port 11 nsew
rlabel metal2 s 278594 279520 278650 280000 6 gpio_dm0[18]
port 12 nsew
rlabel metal2 s 230018 279520 230074 280000 6 gpio_dm0[19]
port 13 nsew
rlabel metal3 s 439520 38632 440000 38752 6 gpio_dm0[1]
port 14 nsew
rlabel metal2 s 181442 279520 181498 280000 6 gpio_dm0[20]
port 15 nsew
rlabel metal2 s 132866 279520 132922 280000 6 gpio_dm0[21]
port 16 nsew
rlabel metal2 s 84290 279520 84346 280000 6 gpio_dm0[22]
port 17 nsew
rlabel metal2 s 35714 279520 35770 280000 6 gpio_dm0[23]
port 18 nsew
rlabel metal3 s 0 272824 480 272944 6 gpio_dm0[24]
port 19 nsew
rlabel metal3 s 0 253240 480 253360 6 gpio_dm0[25]
port 20 nsew
rlabel metal3 s 0 233656 480 233776 6 gpio_dm0[26]
port 21 nsew
rlabel metal3 s 0 214072 480 214192 6 gpio_dm0[27]
port 22 nsew
rlabel metal3 s 0 194488 480 194608 6 gpio_dm0[28]
port 23 nsew
rlabel metal3 s 0 174904 480 175024 6 gpio_dm0[29]
port 24 nsew
rlabel metal3 s 439520 54952 440000 55072 6 gpio_dm0[2]
port 25 nsew
rlabel metal3 s 0 155320 480 155440 6 gpio_dm0[30]
port 26 nsew
rlabel metal3 s 0 135736 480 135856 6 gpio_dm0[31]
port 27 nsew
rlabel metal3 s 0 116152 480 116272 6 gpio_dm0[32]
port 28 nsew
rlabel metal3 s 0 96568 480 96688 6 gpio_dm0[33]
port 29 nsew
rlabel metal3 s 0 76984 480 77104 6 gpio_dm0[34]
port 30 nsew
rlabel metal3 s 0 57400 480 57520 6 gpio_dm0[35]
port 31 nsew
rlabel metal3 s 0 37816 480 37936 6 gpio_dm0[36]
port 32 nsew
rlabel metal3 s 0 18232 480 18352 6 gpio_dm0[37]
port 33 nsew
rlabel metal2 s 21178 0 21234 480 6 gpio_dm0[38]
port 34 nsew
rlabel metal2 s 70858 0 70914 480 6 gpio_dm0[39]
port 35 nsew
rlabel metal3 s 439520 71272 440000 71392 6 gpio_dm0[3]
port 36 nsew
rlabel metal2 s 120538 0 120594 480 6 gpio_dm0[40]
port 37 nsew
rlabel metal2 s 170218 0 170274 480 6 gpio_dm0[41]
port 38 nsew
rlabel metal2 s 219898 0 219954 480 6 gpio_dm0[42]
port 39 nsew
rlabel metal2 s 269578 0 269634 480 6 gpio_dm0[43]
port 40 nsew
rlabel metal3 s 439520 87592 440000 87712 6 gpio_dm0[4]
port 41 nsew
rlabel metal3 s 439520 103912 440000 104032 6 gpio_dm0[5]
port 42 nsew
rlabel metal3 s 439520 120232 440000 120352 6 gpio_dm0[6]
port 43 nsew
rlabel metal3 s 439520 136552 440000 136672 6 gpio_dm0[7]
port 44 nsew
rlabel metal3 s 439520 152872 440000 152992 6 gpio_dm0[8]
port 45 nsew
rlabel metal3 s 439520 169192 440000 169312 6 gpio_dm0[9]
port 46 nsew
rlabel metal3 s 439520 20952 440000 21072 6 gpio_dm1[0]
port 47 nsew
rlabel metal3 s 439520 184152 440000 184272 6 gpio_dm1[10]
port 48 nsew
rlabel metal3 s 439520 200472 440000 200592 6 gpio_dm1[11]
port 49 nsew
rlabel metal3 s 439520 216792 440000 216912 6 gpio_dm1[12]
port 50 nsew
rlabel metal3 s 439520 233112 440000 233232 6 gpio_dm1[13]
port 51 nsew
rlabel metal3 s 439520 249432 440000 249552 6 gpio_dm1[14]
port 52 nsew
rlabel metal2 s 428370 279520 428426 280000 6 gpio_dm1[15]
port 53 nsew
rlabel metal2 s 379794 279520 379850 280000 6 gpio_dm1[16]
port 54 nsew
rlabel metal2 s 331218 279520 331274 280000 6 gpio_dm1[17]
port 55 nsew
rlabel metal2 s 282642 279520 282698 280000 6 gpio_dm1[18]
port 56 nsew
rlabel metal2 s 234066 279520 234122 280000 6 gpio_dm1[19]
port 57 nsew
rlabel metal3 s 439520 37272 440000 37392 6 gpio_dm1[1]
port 58 nsew
rlabel metal2 s 185490 279520 185546 280000 6 gpio_dm1[20]
port 59 nsew
rlabel metal2 s 136914 279520 136970 280000 6 gpio_dm1[21]
port 60 nsew
rlabel metal2 s 88338 279520 88394 280000 6 gpio_dm1[22]
port 61 nsew
rlabel metal2 s 39762 279520 39818 280000 6 gpio_dm1[23]
port 62 nsew
rlabel metal3 s 0 274456 480 274576 6 gpio_dm1[24]
port 63 nsew
rlabel metal3 s 0 254872 480 254992 6 gpio_dm1[25]
port 64 nsew
rlabel metal3 s 0 235288 480 235408 6 gpio_dm1[26]
port 65 nsew
rlabel metal3 s 0 215704 480 215824 6 gpio_dm1[27]
port 66 nsew
rlabel metal3 s 0 196120 480 196240 6 gpio_dm1[28]
port 67 nsew
rlabel metal3 s 0 176536 480 176656 6 gpio_dm1[29]
port 68 nsew
rlabel metal3 s 439520 53592 440000 53712 6 gpio_dm1[2]
port 69 nsew
rlabel metal3 s 0 156952 480 157072 6 gpio_dm1[30]
port 70 nsew
rlabel metal3 s 0 137368 480 137488 6 gpio_dm1[31]
port 71 nsew
rlabel metal3 s 0 117784 480 117904 6 gpio_dm1[32]
port 72 nsew
rlabel metal3 s 0 98200 480 98320 6 gpio_dm1[33]
port 73 nsew
rlabel metal3 s 0 78616 480 78736 6 gpio_dm1[34]
port 74 nsew
rlabel metal3 s 0 59032 480 59152 6 gpio_dm1[35]
port 75 nsew
rlabel metal3 s 0 39448 480 39568 6 gpio_dm1[36]
port 76 nsew
rlabel metal3 s 0 19864 480 19984 6 gpio_dm1[37]
port 77 nsew
rlabel metal2 s 17038 0 17094 480 6 gpio_dm1[38]
port 78 nsew
rlabel metal2 s 66718 0 66774 480 6 gpio_dm1[39]
port 79 nsew
rlabel metal3 s 439520 69912 440000 70032 6 gpio_dm1[3]
port 80 nsew
rlabel metal2 s 116398 0 116454 480 6 gpio_dm1[40]
port 81 nsew
rlabel metal2 s 166078 0 166134 480 6 gpio_dm1[41]
port 82 nsew
rlabel metal2 s 215758 0 215814 480 6 gpio_dm1[42]
port 83 nsew
rlabel metal2 s 265438 0 265494 480 6 gpio_dm1[43]
port 84 nsew
rlabel metal3 s 439520 86232 440000 86352 6 gpio_dm1[4]
port 85 nsew
rlabel metal3 s 439520 102552 440000 102672 6 gpio_dm1[5]
port 86 nsew
rlabel metal3 s 439520 118872 440000 118992 6 gpio_dm1[6]
port 87 nsew
rlabel metal3 s 439520 135192 440000 135312 6 gpio_dm1[7]
port 88 nsew
rlabel metal3 s 439520 151512 440000 151632 6 gpio_dm1[8]
port 89 nsew
rlabel metal3 s 439520 167832 440000 167952 6 gpio_dm1[9]
port 90 nsew
rlabel metal3 s 439520 25032 440000 25152 6 gpio_dm2[0]
port 91 nsew
rlabel metal3 s 439520 188232 440000 188352 6 gpio_dm2[10]
port 92 nsew
rlabel metal3 s 439520 204552 440000 204672 6 gpio_dm2[11]
port 93 nsew
rlabel metal3 s 439520 220872 440000 220992 6 gpio_dm2[12]
port 94 nsew
rlabel metal3 s 439520 237192 440000 237312 6 gpio_dm2[13]
port 95 nsew
rlabel metal3 s 439520 253512 440000 253632 6 gpio_dm2[14]
port 96 nsew
rlabel metal2 s 416226 279520 416282 280000 6 gpio_dm2[15]
port 97 nsew
rlabel metal2 s 367650 279520 367706 280000 6 gpio_dm2[16]
port 98 nsew
rlabel metal2 s 319074 279520 319130 280000 6 gpio_dm2[17]
port 99 nsew
rlabel metal2 s 270498 279520 270554 280000 6 gpio_dm2[18]
port 100 nsew
rlabel metal2 s 221922 279520 221978 280000 6 gpio_dm2[19]
port 101 nsew
rlabel metal3 s 439520 41352 440000 41472 6 gpio_dm2[1]
port 102 nsew
rlabel metal2 s 173346 279520 173402 280000 6 gpio_dm2[20]
port 103 nsew
rlabel metal2 s 124770 279520 124826 280000 6 gpio_dm2[21]
port 104 nsew
rlabel metal2 s 76194 279520 76250 280000 6 gpio_dm2[22]
port 105 nsew
rlabel metal2 s 27618 279520 27674 280000 6 gpio_dm2[23]
port 106 nsew
rlabel metal3 s 0 269560 480 269680 6 gpio_dm2[24]
port 107 nsew
rlabel metal3 s 0 249976 480 250096 6 gpio_dm2[25]
port 108 nsew
rlabel metal3 s 0 230392 480 230512 6 gpio_dm2[26]
port 109 nsew
rlabel metal3 s 0 210808 480 210928 6 gpio_dm2[27]
port 110 nsew
rlabel metal3 s 0 191224 480 191344 6 gpio_dm2[28]
port 111 nsew
rlabel metal3 s 0 171640 480 171760 6 gpio_dm2[29]
port 112 nsew
rlabel metal3 s 439520 57672 440000 57792 6 gpio_dm2[2]
port 113 nsew
rlabel metal3 s 0 152056 480 152176 6 gpio_dm2[30]
port 114 nsew
rlabel metal3 s 0 132472 480 132592 6 gpio_dm2[31]
port 115 nsew
rlabel metal3 s 0 112888 480 113008 6 gpio_dm2[32]
port 116 nsew
rlabel metal3 s 0 93304 480 93424 6 gpio_dm2[33]
port 117 nsew
rlabel metal3 s 0 73720 480 73840 6 gpio_dm2[34]
port 118 nsew
rlabel metal3 s 0 54136 480 54256 6 gpio_dm2[35]
port 119 nsew
rlabel metal3 s 0 34552 480 34672 6 gpio_dm2[36]
port 120 nsew
rlabel metal3 s 0 14968 480 15088 6 gpio_dm2[37]
port 121 nsew
rlabel metal2 s 29458 0 29514 480 6 gpio_dm2[38]
port 122 nsew
rlabel metal2 s 79138 0 79194 480 6 gpio_dm2[39]
port 123 nsew
rlabel metal3 s 439520 73992 440000 74112 6 gpio_dm2[3]
port 124 nsew
rlabel metal2 s 128818 0 128874 480 6 gpio_dm2[40]
port 125 nsew
rlabel metal2 s 178498 0 178554 480 6 gpio_dm2[41]
port 126 nsew
rlabel metal2 s 228178 0 228234 480 6 gpio_dm2[42]
port 127 nsew
rlabel metal2 s 277858 0 277914 480 6 gpio_dm2[43]
port 128 nsew
rlabel metal3 s 439520 90312 440000 90432 6 gpio_dm2[4]
port 129 nsew
rlabel metal3 s 439520 106632 440000 106752 6 gpio_dm2[5]
port 130 nsew
rlabel metal3 s 439520 122952 440000 123072 6 gpio_dm2[6]
port 131 nsew
rlabel metal3 s 439520 139272 440000 139392 6 gpio_dm2[7]
port 132 nsew
rlabel metal3 s 439520 155592 440000 155712 6 gpio_dm2[8]
port 133 nsew
rlabel metal3 s 439520 171912 440000 172032 6 gpio_dm2[9]
port 134 nsew
rlabel metal3 s 439520 29112 440000 29232 6 gpio_ib_mode_sel[0]
port 135 nsew
rlabel metal3 s 439520 192312 440000 192432 6 gpio_ib_mode_sel[10]
port 136 nsew
rlabel metal3 s 439520 208632 440000 208752 6 gpio_ib_mode_sel[11]
port 137 nsew
rlabel metal3 s 439520 224952 440000 225072 6 gpio_ib_mode_sel[12]
port 138 nsew
rlabel metal3 s 439520 241272 440000 241392 6 gpio_ib_mode_sel[13]
port 139 nsew
rlabel metal3 s 439520 257592 440000 257712 6 gpio_ib_mode_sel[14]
port 140 nsew
rlabel metal2 s 404082 279520 404138 280000 6 gpio_ib_mode_sel[15]
port 141 nsew
rlabel metal2 s 355506 279520 355562 280000 6 gpio_ib_mode_sel[16]
port 142 nsew
rlabel metal2 s 306930 279520 306986 280000 6 gpio_ib_mode_sel[17]
port 143 nsew
rlabel metal2 s 258354 279520 258410 280000 6 gpio_ib_mode_sel[18]
port 144 nsew
rlabel metal2 s 209778 279520 209834 280000 6 gpio_ib_mode_sel[19]
port 145 nsew
rlabel metal3 s 439520 45432 440000 45552 6 gpio_ib_mode_sel[1]
port 146 nsew
rlabel metal2 s 161202 279520 161258 280000 6 gpio_ib_mode_sel[20]
port 147 nsew
rlabel metal2 s 112626 279520 112682 280000 6 gpio_ib_mode_sel[21]
port 148 nsew
rlabel metal2 s 64050 279520 64106 280000 6 gpio_ib_mode_sel[22]
port 149 nsew
rlabel metal2 s 15474 279520 15530 280000 6 gpio_ib_mode_sel[23]
port 150 nsew
rlabel metal3 s 0 264664 480 264784 6 gpio_ib_mode_sel[24]
port 151 nsew
rlabel metal3 s 0 245080 480 245200 6 gpio_ib_mode_sel[25]
port 152 nsew
rlabel metal3 s 0 225496 480 225616 6 gpio_ib_mode_sel[26]
port 153 nsew
rlabel metal3 s 0 205912 480 206032 6 gpio_ib_mode_sel[27]
port 154 nsew
rlabel metal3 s 0 186328 480 186448 6 gpio_ib_mode_sel[28]
port 155 nsew
rlabel metal3 s 0 166744 480 166864 6 gpio_ib_mode_sel[29]
port 156 nsew
rlabel metal3 s 439520 61752 440000 61872 6 gpio_ib_mode_sel[2]
port 157 nsew
rlabel metal3 s 0 147160 480 147280 6 gpio_ib_mode_sel[30]
port 158 nsew
rlabel metal3 s 0 127576 480 127696 6 gpio_ib_mode_sel[31]
port 159 nsew
rlabel metal3 s 0 107992 480 108112 6 gpio_ib_mode_sel[32]
port 160 nsew
rlabel metal3 s 0 88408 480 88528 6 gpio_ib_mode_sel[33]
port 161 nsew
rlabel metal3 s 0 68824 480 68944 6 gpio_ib_mode_sel[34]
port 162 nsew
rlabel metal3 s 0 49240 480 49360 6 gpio_ib_mode_sel[35]
port 163 nsew
rlabel metal3 s 0 29656 480 29776 6 gpio_ib_mode_sel[36]
port 164 nsew
rlabel metal3 s 0 10072 480 10192 6 gpio_ib_mode_sel[37]
port 165 nsew
rlabel metal2 s 41878 0 41934 480 6 gpio_ib_mode_sel[38]
port 166 nsew
rlabel metal2 s 91558 0 91614 480 6 gpio_ib_mode_sel[39]
port 167 nsew
rlabel metal3 s 439520 78072 440000 78192 6 gpio_ib_mode_sel[3]
port 168 nsew
rlabel metal2 s 141238 0 141294 480 6 gpio_ib_mode_sel[40]
port 169 nsew
rlabel metal2 s 190918 0 190974 480 6 gpio_ib_mode_sel[41]
port 170 nsew
rlabel metal2 s 240598 0 240654 480 6 gpio_ib_mode_sel[42]
port 171 nsew
rlabel metal2 s 290278 0 290334 480 6 gpio_ib_mode_sel[43]
port 172 nsew
rlabel metal3 s 439520 94392 440000 94512 6 gpio_ib_mode_sel[4]
port 173 nsew
rlabel metal3 s 439520 110712 440000 110832 6 gpio_ib_mode_sel[5]
port 174 nsew
rlabel metal3 s 439520 127032 440000 127152 6 gpio_ib_mode_sel[6]
port 175 nsew
rlabel metal3 s 439520 143352 440000 143472 6 gpio_ib_mode_sel[7]
port 176 nsew
rlabel metal3 s 439520 159672 440000 159792 6 gpio_ib_mode_sel[8]
port 177 nsew
rlabel metal3 s 439520 175992 440000 176112 6 gpio_ib_mode_sel[9]
port 178 nsew
rlabel metal3 s 439520 23672 440000 23792 6 gpio_ieb[0]
port 179 nsew
rlabel metal3 s 439520 186872 440000 186992 6 gpio_ieb[10]
port 180 nsew
rlabel metal3 s 439520 203192 440000 203312 6 gpio_ieb[11]
port 181 nsew
rlabel metal3 s 439520 219512 440000 219632 6 gpio_ieb[12]
port 182 nsew
rlabel metal3 s 439520 235832 440000 235952 6 gpio_ieb[13]
port 183 nsew
rlabel metal3 s 439520 252152 440000 252272 6 gpio_ieb[14]
port 184 nsew
rlabel metal2 s 420274 279520 420330 280000 6 gpio_ieb[15]
port 185 nsew
rlabel metal2 s 371698 279520 371754 280000 6 gpio_ieb[16]
port 186 nsew
rlabel metal2 s 323122 279520 323178 280000 6 gpio_ieb[17]
port 187 nsew
rlabel metal2 s 274546 279520 274602 280000 6 gpio_ieb[18]
port 188 nsew
rlabel metal2 s 225970 279520 226026 280000 6 gpio_ieb[19]
port 189 nsew
rlabel metal3 s 439520 39992 440000 40112 6 gpio_ieb[1]
port 190 nsew
rlabel metal2 s 177394 279520 177450 280000 6 gpio_ieb[20]
port 191 nsew
rlabel metal2 s 128818 279520 128874 280000 6 gpio_ieb[21]
port 192 nsew
rlabel metal2 s 80242 279520 80298 280000 6 gpio_ieb[22]
port 193 nsew
rlabel metal2 s 31666 279520 31722 280000 6 gpio_ieb[23]
port 194 nsew
rlabel metal3 s 0 271192 480 271312 6 gpio_ieb[24]
port 195 nsew
rlabel metal3 s 0 251608 480 251728 6 gpio_ieb[25]
port 196 nsew
rlabel metal3 s 0 232024 480 232144 6 gpio_ieb[26]
port 197 nsew
rlabel metal3 s 0 212440 480 212560 6 gpio_ieb[27]
port 198 nsew
rlabel metal3 s 0 192856 480 192976 6 gpio_ieb[28]
port 199 nsew
rlabel metal3 s 0 173272 480 173392 6 gpio_ieb[29]
port 200 nsew
rlabel metal3 s 439520 56312 440000 56432 6 gpio_ieb[2]
port 201 nsew
rlabel metal3 s 0 153688 480 153808 6 gpio_ieb[30]
port 202 nsew
rlabel metal3 s 0 134104 480 134224 6 gpio_ieb[31]
port 203 nsew
rlabel metal3 s 0 114520 480 114640 6 gpio_ieb[32]
port 204 nsew
rlabel metal3 s 0 94936 480 95056 6 gpio_ieb[33]
port 205 nsew
rlabel metal3 s 0 75352 480 75472 6 gpio_ieb[34]
port 206 nsew
rlabel metal3 s 0 55768 480 55888 6 gpio_ieb[35]
port 207 nsew
rlabel metal3 s 0 36184 480 36304 6 gpio_ieb[36]
port 208 nsew
rlabel metal3 s 0 16600 480 16720 6 gpio_ieb[37]
port 209 nsew
rlabel metal2 s 25318 0 25374 480 6 gpio_ieb[38]
port 210 nsew
rlabel metal2 s 74998 0 75054 480 6 gpio_ieb[39]
port 211 nsew
rlabel metal3 s 439520 72632 440000 72752 6 gpio_ieb[3]
port 212 nsew
rlabel metal2 s 124678 0 124734 480 6 gpio_ieb[40]
port 213 nsew
rlabel metal2 s 174358 0 174414 480 6 gpio_ieb[41]
port 214 nsew
rlabel metal2 s 224038 0 224094 480 6 gpio_ieb[42]
port 215 nsew
rlabel metal2 s 273718 0 273774 480 6 gpio_ieb[43]
port 216 nsew
rlabel metal3 s 439520 88952 440000 89072 6 gpio_ieb[4]
port 217 nsew
rlabel metal3 s 439520 105272 440000 105392 6 gpio_ieb[5]
port 218 nsew
rlabel metal3 s 439520 121592 440000 121712 6 gpio_ieb[6]
port 219 nsew
rlabel metal3 s 439520 137912 440000 138032 6 gpio_ieb[7]
port 220 nsew
rlabel metal3 s 439520 154232 440000 154352 6 gpio_ieb[8]
port 221 nsew
rlabel metal3 s 439520 170552 440000 170672 6 gpio_ieb[9]
port 222 nsew
rlabel metal3 s 439520 18232 440000 18352 6 gpio_in[0]
port 223 nsew
rlabel metal3 s 439520 181432 440000 181552 6 gpio_in[10]
port 224 nsew
rlabel metal3 s 439520 197752 440000 197872 6 gpio_in[11]
port 225 nsew
rlabel metal3 s 439520 214072 440000 214192 6 gpio_in[12]
port 226 nsew
rlabel metal3 s 439520 230392 440000 230512 6 gpio_in[13]
port 227 nsew
rlabel metal3 s 439520 246712 440000 246832 6 gpio_in[14]
port 228 nsew
rlabel metal2 s 436466 279520 436522 280000 6 gpio_in[15]
port 229 nsew
rlabel metal2 s 387890 279520 387946 280000 6 gpio_in[16]
port 230 nsew
rlabel metal2 s 339314 279520 339370 280000 6 gpio_in[17]
port 231 nsew
rlabel metal2 s 290738 279520 290794 280000 6 gpio_in[18]
port 232 nsew
rlabel metal2 s 242162 279520 242218 280000 6 gpio_in[19]
port 233 nsew
rlabel metal3 s 439520 34552 440000 34672 6 gpio_in[1]
port 234 nsew
rlabel metal2 s 193586 279520 193642 280000 6 gpio_in[20]
port 235 nsew
rlabel metal2 s 145010 279520 145066 280000 6 gpio_in[21]
port 236 nsew
rlabel metal2 s 96434 279520 96490 280000 6 gpio_in[22]
port 237 nsew
rlabel metal2 s 47858 279520 47914 280000 6 gpio_in[23]
port 238 nsew
rlabel metal3 s 0 277720 480 277840 6 gpio_in[24]
port 239 nsew
rlabel metal3 s 0 258136 480 258256 6 gpio_in[25]
port 240 nsew
rlabel metal3 s 0 238552 480 238672 6 gpio_in[26]
port 241 nsew
rlabel metal3 s 0 218968 480 219088 6 gpio_in[27]
port 242 nsew
rlabel metal3 s 0 199384 480 199504 6 gpio_in[28]
port 243 nsew
rlabel metal3 s 0 179800 480 179920 6 gpio_in[29]
port 244 nsew
rlabel metal3 s 439520 50872 440000 50992 6 gpio_in[2]
port 245 nsew
rlabel metal3 s 0 160216 480 160336 6 gpio_in[30]
port 246 nsew
rlabel metal3 s 0 140632 480 140752 6 gpio_in[31]
port 247 nsew
rlabel metal3 s 0 121048 480 121168 6 gpio_in[32]
port 248 nsew
rlabel metal3 s 0 101464 480 101584 6 gpio_in[33]
port 249 nsew
rlabel metal3 s 0 81880 480 82000 6 gpio_in[34]
port 250 nsew
rlabel metal3 s 0 62296 480 62416 6 gpio_in[35]
port 251 nsew
rlabel metal3 s 0 42712 480 42832 6 gpio_in[36]
port 252 nsew
rlabel metal3 s 0 23128 480 23248 6 gpio_in[37]
port 253 nsew
rlabel metal2 s 8758 0 8814 480 6 gpio_in[38]
port 254 nsew
rlabel metal2 s 58438 0 58494 480 6 gpio_in[39]
port 255 nsew
rlabel metal3 s 439520 67192 440000 67312 6 gpio_in[3]
port 256 nsew
rlabel metal2 s 108118 0 108174 480 6 gpio_in[40]
port 257 nsew
rlabel metal2 s 157798 0 157854 480 6 gpio_in[41]
port 258 nsew
rlabel metal2 s 207478 0 207534 480 6 gpio_in[42]
port 259 nsew
rlabel metal2 s 257158 0 257214 480 6 gpio_in[43]
port 260 nsew
rlabel metal3 s 439520 83512 440000 83632 6 gpio_in[4]
port 261 nsew
rlabel metal3 s 439520 99832 440000 99952 6 gpio_in[5]
port 262 nsew
rlabel metal3 s 439520 116152 440000 116272 6 gpio_in[6]
port 263 nsew
rlabel metal3 s 439520 132472 440000 132592 6 gpio_in[7]
port 264 nsew
rlabel metal3 s 439520 148792 440000 148912 6 gpio_in[8]
port 265 nsew
rlabel metal3 s 439520 165112 440000 165232 6 gpio_in[9]
port 266 nsew
rlabel metal3 s 439520 31832 440000 31952 6 gpio_loopback_one[0]
port 267 nsew
rlabel metal3 s 439520 195032 440000 195152 6 gpio_loopback_one[10]
port 268 nsew
rlabel metal3 s 439520 211352 440000 211472 6 gpio_loopback_one[11]
port 269 nsew
rlabel metal3 s 439520 227672 440000 227792 6 gpio_loopback_one[12]
port 270 nsew
rlabel metal3 s 439520 243992 440000 244112 6 gpio_loopback_one[13]
port 271 nsew
rlabel metal3 s 439520 260312 440000 260432 6 gpio_loopback_one[14]
port 272 nsew
rlabel metal2 s 395986 279520 396042 280000 6 gpio_loopback_one[15]
port 273 nsew
rlabel metal2 s 347410 279520 347466 280000 6 gpio_loopback_one[16]
port 274 nsew
rlabel metal2 s 298834 279520 298890 280000 6 gpio_loopback_one[17]
port 275 nsew
rlabel metal2 s 250258 279520 250314 280000 6 gpio_loopback_one[18]
port 276 nsew
rlabel metal2 s 201682 279520 201738 280000 6 gpio_loopback_one[19]
port 277 nsew
rlabel metal3 s 439520 48152 440000 48272 6 gpio_loopback_one[1]
port 278 nsew
rlabel metal2 s 153106 279520 153162 280000 6 gpio_loopback_one[20]
port 279 nsew
rlabel metal2 s 104530 279520 104586 280000 6 gpio_loopback_one[21]
port 280 nsew
rlabel metal2 s 55954 279520 56010 280000 6 gpio_loopback_one[22]
port 281 nsew
rlabel metal2 s 7378 279520 7434 280000 6 gpio_loopback_one[23]
port 282 nsew
rlabel metal3 s 0 261400 480 261520 6 gpio_loopback_one[24]
port 283 nsew
rlabel metal3 s 0 241816 480 241936 6 gpio_loopback_one[25]
port 284 nsew
rlabel metal3 s 0 222232 480 222352 6 gpio_loopback_one[26]
port 285 nsew
rlabel metal3 s 0 202648 480 202768 6 gpio_loopback_one[27]
port 286 nsew
rlabel metal3 s 0 183064 480 183184 6 gpio_loopback_one[28]
port 287 nsew
rlabel metal3 s 0 163480 480 163600 6 gpio_loopback_one[29]
port 288 nsew
rlabel metal3 s 439520 64472 440000 64592 6 gpio_loopback_one[2]
port 289 nsew
rlabel metal3 s 0 143896 480 144016 6 gpio_loopback_one[30]
port 290 nsew
rlabel metal3 s 0 124312 480 124432 6 gpio_loopback_one[31]
port 291 nsew
rlabel metal3 s 0 104728 480 104848 6 gpio_loopback_one[32]
port 292 nsew
rlabel metal3 s 0 85144 480 85264 6 gpio_loopback_one[33]
port 293 nsew
rlabel metal3 s 0 65560 480 65680 6 gpio_loopback_one[34]
port 294 nsew
rlabel metal3 s 0 45976 480 46096 6 gpio_loopback_one[35]
port 295 nsew
rlabel metal3 s 0 26392 480 26512 6 gpio_loopback_one[36]
port 296 nsew
rlabel metal3 s 0 6808 480 6928 6 gpio_loopback_one[37]
port 297 nsew
rlabel metal2 s 50158 0 50214 480 6 gpio_loopback_one[38]
port 298 nsew
rlabel metal2 s 99838 0 99894 480 6 gpio_loopback_one[39]
port 299 nsew
rlabel metal3 s 439520 80792 440000 80912 6 gpio_loopback_one[3]
port 300 nsew
rlabel metal2 s 149518 0 149574 480 6 gpio_loopback_one[40]
port 301 nsew
rlabel metal2 s 199198 0 199254 480 6 gpio_loopback_one[41]
port 302 nsew
rlabel metal2 s 248878 0 248934 480 6 gpio_loopback_one[42]
port 303 nsew
rlabel metal2 s 298558 0 298614 480 6 gpio_loopback_one[43]
port 304 nsew
rlabel metal3 s 439520 97112 440000 97232 6 gpio_loopback_one[4]
port 305 nsew
rlabel metal3 s 439520 113432 440000 113552 6 gpio_loopback_one[5]
port 306 nsew
rlabel metal3 s 439520 129752 440000 129872 6 gpio_loopback_one[6]
port 307 nsew
rlabel metal3 s 439520 146072 440000 146192 6 gpio_loopback_one[7]
port 308 nsew
rlabel metal3 s 439520 162392 440000 162512 6 gpio_loopback_one[8]
port 309 nsew
rlabel metal3 s 439520 178712 440000 178832 6 gpio_loopback_one[9]
port 310 nsew
rlabel metal3 s 439520 33192 440000 33312 6 gpio_loopback_zero[0]
port 311 nsew
rlabel metal3 s 439520 196392 440000 196512 6 gpio_loopback_zero[10]
port 312 nsew
rlabel metal3 s 439520 212712 440000 212832 6 gpio_loopback_zero[11]
port 313 nsew
rlabel metal3 s 439520 229032 440000 229152 6 gpio_loopback_zero[12]
port 314 nsew
rlabel metal3 s 439520 245352 440000 245472 6 gpio_loopback_zero[13]
port 315 nsew
rlabel metal3 s 439520 261672 440000 261792 6 gpio_loopback_zero[14]
port 316 nsew
rlabel metal2 s 391938 279520 391994 280000 6 gpio_loopback_zero[15]
port 317 nsew
rlabel metal2 s 343362 279520 343418 280000 6 gpio_loopback_zero[16]
port 318 nsew
rlabel metal2 s 294786 279520 294842 280000 6 gpio_loopback_zero[17]
port 319 nsew
rlabel metal2 s 246210 279520 246266 280000 6 gpio_loopback_zero[18]
port 320 nsew
rlabel metal2 s 197634 279520 197690 280000 6 gpio_loopback_zero[19]
port 321 nsew
rlabel metal3 s 439520 49512 440000 49632 6 gpio_loopback_zero[1]
port 322 nsew
rlabel metal2 s 149058 279520 149114 280000 6 gpio_loopback_zero[20]
port 323 nsew
rlabel metal2 s 100482 279520 100538 280000 6 gpio_loopback_zero[21]
port 324 nsew
rlabel metal2 s 51906 279520 51962 280000 6 gpio_loopback_zero[22]
port 325 nsew
rlabel metal2 s 3330 279520 3386 280000 6 gpio_loopback_zero[23]
port 326 nsew
rlabel metal3 s 0 259768 480 259888 6 gpio_loopback_zero[24]
port 327 nsew
rlabel metal3 s 0 240184 480 240304 6 gpio_loopback_zero[25]
port 328 nsew
rlabel metal3 s 0 220600 480 220720 6 gpio_loopback_zero[26]
port 329 nsew
rlabel metal3 s 0 201016 480 201136 6 gpio_loopback_zero[27]
port 330 nsew
rlabel metal3 s 0 181432 480 181552 6 gpio_loopback_zero[28]
port 331 nsew
rlabel metal3 s 0 161848 480 161968 6 gpio_loopback_zero[29]
port 332 nsew
rlabel metal3 s 439520 65832 440000 65952 6 gpio_loopback_zero[2]
port 333 nsew
rlabel metal3 s 0 142264 480 142384 6 gpio_loopback_zero[30]
port 334 nsew
rlabel metal3 s 0 122680 480 122800 6 gpio_loopback_zero[31]
port 335 nsew
rlabel metal3 s 0 103096 480 103216 6 gpio_loopback_zero[32]
port 336 nsew
rlabel metal3 s 0 83512 480 83632 6 gpio_loopback_zero[33]
port 337 nsew
rlabel metal3 s 0 63928 480 64048 6 gpio_loopback_zero[34]
port 338 nsew
rlabel metal3 s 0 44344 480 44464 6 gpio_loopback_zero[35]
port 339 nsew
rlabel metal3 s 0 24760 480 24880 6 gpio_loopback_zero[36]
port 340 nsew
rlabel metal3 s 0 5176 480 5296 6 gpio_loopback_zero[37]
port 341 nsew
rlabel metal2 s 54298 0 54354 480 6 gpio_loopback_zero[38]
port 342 nsew
rlabel metal2 s 103978 0 104034 480 6 gpio_loopback_zero[39]
port 343 nsew
rlabel metal3 s 439520 82152 440000 82272 6 gpio_loopback_zero[3]
port 344 nsew
rlabel metal2 s 153658 0 153714 480 6 gpio_loopback_zero[40]
port 345 nsew
rlabel metal2 s 203338 0 203394 480 6 gpio_loopback_zero[41]
port 346 nsew
rlabel metal2 s 253018 0 253074 480 6 gpio_loopback_zero[42]
port 347 nsew
rlabel metal2 s 302698 0 302754 480 6 gpio_loopback_zero[43]
port 348 nsew
rlabel metal3 s 439520 98472 440000 98592 6 gpio_loopback_zero[4]
port 349 nsew
rlabel metal3 s 439520 114792 440000 114912 6 gpio_loopback_zero[5]
port 350 nsew
rlabel metal3 s 439520 131112 440000 131232 6 gpio_loopback_zero[6]
port 351 nsew
rlabel metal3 s 439520 147432 440000 147552 6 gpio_loopback_zero[7]
port 352 nsew
rlabel metal3 s 439520 163752 440000 163872 6 gpio_loopback_zero[8]
port 353 nsew
rlabel metal3 s 439520 180072 440000 180192 6 gpio_loopback_zero[9]
port 354 nsew
rlabel metal3 s 439520 30472 440000 30592 6 gpio_oeb[0]
port 355 nsew
rlabel metal3 s 439520 193672 440000 193792 6 gpio_oeb[10]
port 356 nsew
rlabel metal3 s 439520 209992 440000 210112 6 gpio_oeb[11]
port 357 nsew
rlabel metal3 s 439520 226312 440000 226432 6 gpio_oeb[12]
port 358 nsew
rlabel metal3 s 439520 242632 440000 242752 6 gpio_oeb[13]
port 359 nsew
rlabel metal3 s 439520 258952 440000 259072 6 gpio_oeb[14]
port 360 nsew
rlabel metal2 s 400034 279520 400090 280000 6 gpio_oeb[15]
port 361 nsew
rlabel metal2 s 351458 279520 351514 280000 6 gpio_oeb[16]
port 362 nsew
rlabel metal2 s 302882 279520 302938 280000 6 gpio_oeb[17]
port 363 nsew
rlabel metal2 s 254306 279520 254362 280000 6 gpio_oeb[18]
port 364 nsew
rlabel metal2 s 205730 279520 205786 280000 6 gpio_oeb[19]
port 365 nsew
rlabel metal3 s 439520 46792 440000 46912 6 gpio_oeb[1]
port 366 nsew
rlabel metal2 s 157154 279520 157210 280000 6 gpio_oeb[20]
port 367 nsew
rlabel metal2 s 108578 279520 108634 280000 6 gpio_oeb[21]
port 368 nsew
rlabel metal2 s 60002 279520 60058 280000 6 gpio_oeb[22]
port 369 nsew
rlabel metal2 s 11426 279520 11482 280000 6 gpio_oeb[23]
port 370 nsew
rlabel metal3 s 0 263032 480 263152 6 gpio_oeb[24]
port 371 nsew
rlabel metal3 s 0 243448 480 243568 6 gpio_oeb[25]
port 372 nsew
rlabel metal3 s 0 223864 480 223984 6 gpio_oeb[26]
port 373 nsew
rlabel metal3 s 0 204280 480 204400 6 gpio_oeb[27]
port 374 nsew
rlabel metal3 s 0 184696 480 184816 6 gpio_oeb[28]
port 375 nsew
rlabel metal3 s 0 165112 480 165232 6 gpio_oeb[29]
port 376 nsew
rlabel metal3 s 439520 63112 440000 63232 6 gpio_oeb[2]
port 377 nsew
rlabel metal3 s 0 145528 480 145648 6 gpio_oeb[30]
port 378 nsew
rlabel metal3 s 0 125944 480 126064 6 gpio_oeb[31]
port 379 nsew
rlabel metal3 s 0 106360 480 106480 6 gpio_oeb[32]
port 380 nsew
rlabel metal3 s 0 86776 480 86896 6 gpio_oeb[33]
port 381 nsew
rlabel metal3 s 0 67192 480 67312 6 gpio_oeb[34]
port 382 nsew
rlabel metal3 s 0 47608 480 47728 6 gpio_oeb[35]
port 383 nsew
rlabel metal3 s 0 28024 480 28144 6 gpio_oeb[36]
port 384 nsew
rlabel metal3 s 0 8440 480 8560 6 gpio_oeb[37]
port 385 nsew
rlabel metal2 s 46018 0 46074 480 6 gpio_oeb[38]
port 386 nsew
rlabel metal2 s 95698 0 95754 480 6 gpio_oeb[39]
port 387 nsew
rlabel metal3 s 439520 79432 440000 79552 6 gpio_oeb[3]
port 388 nsew
rlabel metal2 s 145378 0 145434 480 6 gpio_oeb[40]
port 389 nsew
rlabel metal2 s 195058 0 195114 480 6 gpio_oeb[41]
port 390 nsew
rlabel metal2 s 244738 0 244794 480 6 gpio_oeb[42]
port 391 nsew
rlabel metal2 s 294418 0 294474 480 6 gpio_oeb[43]
port 392 nsew
rlabel metal3 s 439520 95752 440000 95872 6 gpio_oeb[4]
port 393 nsew
rlabel metal3 s 439520 112072 440000 112192 6 gpio_oeb[5]
port 394 nsew
rlabel metal3 s 439520 128392 440000 128512 6 gpio_oeb[6]
port 395 nsew
rlabel metal3 s 439520 144712 440000 144832 6 gpio_oeb[7]
port 396 nsew
rlabel metal3 s 439520 161032 440000 161152 6 gpio_oeb[8]
port 397 nsew
rlabel metal3 s 439520 177352 440000 177472 6 gpio_oeb[9]
port 398 nsew
rlabel metal3 s 439520 26392 440000 26512 6 gpio_out[0]
port 399 nsew
rlabel metal3 s 439520 189592 440000 189712 6 gpio_out[10]
port 400 nsew
rlabel metal3 s 439520 205912 440000 206032 6 gpio_out[11]
port 401 nsew
rlabel metal3 s 439520 222232 440000 222352 6 gpio_out[12]
port 402 nsew
rlabel metal3 s 439520 238552 440000 238672 6 gpio_out[13]
port 403 nsew
rlabel metal3 s 439520 254872 440000 254992 6 gpio_out[14]
port 404 nsew
rlabel metal2 s 412178 279520 412234 280000 6 gpio_out[15]
port 405 nsew
rlabel metal2 s 363602 279520 363658 280000 6 gpio_out[16]
port 406 nsew
rlabel metal2 s 315026 279520 315082 280000 6 gpio_out[17]
port 407 nsew
rlabel metal2 s 266450 279520 266506 280000 6 gpio_out[18]
port 408 nsew
rlabel metal2 s 217874 279520 217930 280000 6 gpio_out[19]
port 409 nsew
rlabel metal3 s 439520 42712 440000 42832 6 gpio_out[1]
port 410 nsew
rlabel metal2 s 169298 279520 169354 280000 6 gpio_out[20]
port 411 nsew
rlabel metal2 s 120722 279520 120778 280000 6 gpio_out[21]
port 412 nsew
rlabel metal2 s 72146 279520 72202 280000 6 gpio_out[22]
port 413 nsew
rlabel metal2 s 23570 279520 23626 280000 6 gpio_out[23]
port 414 nsew
rlabel metal3 s 0 267928 480 268048 6 gpio_out[24]
port 415 nsew
rlabel metal3 s 0 248344 480 248464 6 gpio_out[25]
port 416 nsew
rlabel metal3 s 0 228760 480 228880 6 gpio_out[26]
port 417 nsew
rlabel metal3 s 0 209176 480 209296 6 gpio_out[27]
port 418 nsew
rlabel metal3 s 0 189592 480 189712 6 gpio_out[28]
port 419 nsew
rlabel metal3 s 0 170008 480 170128 6 gpio_out[29]
port 420 nsew
rlabel metal3 s 439520 59032 440000 59152 6 gpio_out[2]
port 421 nsew
rlabel metal3 s 0 150424 480 150544 6 gpio_out[30]
port 422 nsew
rlabel metal3 s 0 130840 480 130960 6 gpio_out[31]
port 423 nsew
rlabel metal3 s 0 111256 480 111376 6 gpio_out[32]
port 424 nsew
rlabel metal3 s 0 91672 480 91792 6 gpio_out[33]
port 425 nsew
rlabel metal3 s 0 72088 480 72208 6 gpio_out[34]
port 426 nsew
rlabel metal3 s 0 52504 480 52624 6 gpio_out[35]
port 427 nsew
rlabel metal3 s 0 32920 480 33040 6 gpio_out[36]
port 428 nsew
rlabel metal3 s 0 13336 480 13456 6 gpio_out[37]
port 429 nsew
rlabel metal2 s 33598 0 33654 480 6 gpio_out[38]
port 430 nsew
rlabel metal2 s 83278 0 83334 480 6 gpio_out[39]
port 431 nsew
rlabel metal3 s 439520 75352 440000 75472 6 gpio_out[3]
port 432 nsew
rlabel metal2 s 132958 0 133014 480 6 gpio_out[40]
port 433 nsew
rlabel metal2 s 182638 0 182694 480 6 gpio_out[41]
port 434 nsew
rlabel metal2 s 232318 0 232374 480 6 gpio_out[42]
port 435 nsew
rlabel metal2 s 281998 0 282054 480 6 gpio_out[43]
port 436 nsew
rlabel metal3 s 439520 91672 440000 91792 6 gpio_out[4]
port 437 nsew
rlabel metal3 s 439520 107992 440000 108112 6 gpio_out[5]
port 438 nsew
rlabel metal3 s 439520 124312 440000 124432 6 gpio_out[6]
port 439 nsew
rlabel metal3 s 439520 140632 440000 140752 6 gpio_out[7]
port 440 nsew
rlabel metal3 s 439520 156952 440000 157072 6 gpio_out[8]
port 441 nsew
rlabel metal3 s 439520 173272 440000 173392 6 gpio_out[9]
port 442 nsew
rlabel metal3 s 439520 19592 440000 19712 6 gpio_slow_sel[0]
port 443 nsew
rlabel metal3 s 439520 182792 440000 182912 6 gpio_slow_sel[10]
port 444 nsew
rlabel metal3 s 439520 199112 440000 199232 6 gpio_slow_sel[11]
port 445 nsew
rlabel metal3 s 439520 215432 440000 215552 6 gpio_slow_sel[12]
port 446 nsew
rlabel metal3 s 439520 231752 440000 231872 6 gpio_slow_sel[13]
port 447 nsew
rlabel metal3 s 439520 248072 440000 248192 6 gpio_slow_sel[14]
port 448 nsew
rlabel metal2 s 432418 279520 432474 280000 6 gpio_slow_sel[15]
port 449 nsew
rlabel metal2 s 383842 279520 383898 280000 6 gpio_slow_sel[16]
port 450 nsew
rlabel metal2 s 335266 279520 335322 280000 6 gpio_slow_sel[17]
port 451 nsew
rlabel metal2 s 286690 279520 286746 280000 6 gpio_slow_sel[18]
port 452 nsew
rlabel metal2 s 238114 279520 238170 280000 6 gpio_slow_sel[19]
port 453 nsew
rlabel metal3 s 439520 35912 440000 36032 6 gpio_slow_sel[1]
port 454 nsew
rlabel metal2 s 189538 279520 189594 280000 6 gpio_slow_sel[20]
port 455 nsew
rlabel metal2 s 140962 279520 141018 280000 6 gpio_slow_sel[21]
port 456 nsew
rlabel metal2 s 92386 279520 92442 280000 6 gpio_slow_sel[22]
port 457 nsew
rlabel metal2 s 43810 279520 43866 280000 6 gpio_slow_sel[23]
port 458 nsew
rlabel metal3 s 0 276088 480 276208 6 gpio_slow_sel[24]
port 459 nsew
rlabel metal3 s 0 256504 480 256624 6 gpio_slow_sel[25]
port 460 nsew
rlabel metal3 s 0 236920 480 237040 6 gpio_slow_sel[26]
port 461 nsew
rlabel metal3 s 0 217336 480 217456 6 gpio_slow_sel[27]
port 462 nsew
rlabel metal3 s 0 197752 480 197872 6 gpio_slow_sel[28]
port 463 nsew
rlabel metal3 s 0 178168 480 178288 6 gpio_slow_sel[29]
port 464 nsew
rlabel metal3 s 439520 52232 440000 52352 6 gpio_slow_sel[2]
port 465 nsew
rlabel metal3 s 0 158584 480 158704 6 gpio_slow_sel[30]
port 466 nsew
rlabel metal3 s 0 139000 480 139120 6 gpio_slow_sel[31]
port 467 nsew
rlabel metal3 s 0 119416 480 119536 6 gpio_slow_sel[32]
port 468 nsew
rlabel metal3 s 0 99832 480 99952 6 gpio_slow_sel[33]
port 469 nsew
rlabel metal3 s 0 80248 480 80368 6 gpio_slow_sel[34]
port 470 nsew
rlabel metal3 s 0 60664 480 60784 6 gpio_slow_sel[35]
port 471 nsew
rlabel metal3 s 0 41080 480 41200 6 gpio_slow_sel[36]
port 472 nsew
rlabel metal3 s 0 21496 480 21616 6 gpio_slow_sel[37]
port 473 nsew
rlabel metal2 s 12898 0 12954 480 6 gpio_slow_sel[38]
port 474 nsew
rlabel metal2 s 62578 0 62634 480 6 gpio_slow_sel[39]
port 475 nsew
rlabel metal3 s 439520 68552 440000 68672 6 gpio_slow_sel[3]
port 476 nsew
rlabel metal2 s 112258 0 112314 480 6 gpio_slow_sel[40]
port 477 nsew
rlabel metal2 s 161938 0 161994 480 6 gpio_slow_sel[41]
port 478 nsew
rlabel metal2 s 211618 0 211674 480 6 gpio_slow_sel[42]
port 479 nsew
rlabel metal2 s 261298 0 261354 480 6 gpio_slow_sel[43]
port 480 nsew
rlabel metal3 s 439520 84872 440000 84992 6 gpio_slow_sel[4]
port 481 nsew
rlabel metal3 s 439520 101192 440000 101312 6 gpio_slow_sel[5]
port 482 nsew
rlabel metal3 s 439520 117512 440000 117632 6 gpio_slow_sel[6]
port 483 nsew
rlabel metal3 s 439520 133832 440000 133952 6 gpio_slow_sel[7]
port 484 nsew
rlabel metal3 s 439520 150152 440000 150272 6 gpio_slow_sel[8]
port 485 nsew
rlabel metal3 s 439520 166472 440000 166592 6 gpio_slow_sel[9]
port 486 nsew
rlabel metal3 s 439520 27752 440000 27872 6 gpio_vtrip_sel[0]
port 487 nsew
rlabel metal3 s 439520 190952 440000 191072 6 gpio_vtrip_sel[10]
port 488 nsew
rlabel metal3 s 439520 207272 440000 207392 6 gpio_vtrip_sel[11]
port 489 nsew
rlabel metal3 s 439520 223592 440000 223712 6 gpio_vtrip_sel[12]
port 490 nsew
rlabel metal3 s 439520 239912 440000 240032 6 gpio_vtrip_sel[13]
port 491 nsew
rlabel metal3 s 439520 256232 440000 256352 6 gpio_vtrip_sel[14]
port 492 nsew
rlabel metal2 s 408130 279520 408186 280000 6 gpio_vtrip_sel[15]
port 493 nsew
rlabel metal2 s 359554 279520 359610 280000 6 gpio_vtrip_sel[16]
port 494 nsew
rlabel metal2 s 310978 279520 311034 280000 6 gpio_vtrip_sel[17]
port 495 nsew
rlabel metal2 s 262402 279520 262458 280000 6 gpio_vtrip_sel[18]
port 496 nsew
rlabel metal2 s 213826 279520 213882 280000 6 gpio_vtrip_sel[19]
port 497 nsew
rlabel metal3 s 439520 44072 440000 44192 6 gpio_vtrip_sel[1]
port 498 nsew
rlabel metal2 s 165250 279520 165306 280000 6 gpio_vtrip_sel[20]
port 499 nsew
rlabel metal2 s 116674 279520 116730 280000 6 gpio_vtrip_sel[21]
port 500 nsew
rlabel metal2 s 68098 279520 68154 280000 6 gpio_vtrip_sel[22]
port 501 nsew
rlabel metal2 s 19522 279520 19578 280000 6 gpio_vtrip_sel[23]
port 502 nsew
rlabel metal3 s 0 266296 480 266416 6 gpio_vtrip_sel[24]
port 503 nsew
rlabel metal3 s 0 246712 480 246832 6 gpio_vtrip_sel[25]
port 504 nsew
rlabel metal3 s 0 227128 480 227248 6 gpio_vtrip_sel[26]
port 505 nsew
rlabel metal3 s 0 207544 480 207664 6 gpio_vtrip_sel[27]
port 506 nsew
rlabel metal3 s 0 187960 480 188080 6 gpio_vtrip_sel[28]
port 507 nsew
rlabel metal3 s 0 168376 480 168496 6 gpio_vtrip_sel[29]
port 508 nsew
rlabel metal3 s 439520 60392 440000 60512 6 gpio_vtrip_sel[2]
port 509 nsew
rlabel metal3 s 0 148792 480 148912 6 gpio_vtrip_sel[30]
port 510 nsew
rlabel metal3 s 0 129208 480 129328 6 gpio_vtrip_sel[31]
port 511 nsew
rlabel metal3 s 0 109624 480 109744 6 gpio_vtrip_sel[32]
port 512 nsew
rlabel metal3 s 0 90040 480 90160 6 gpio_vtrip_sel[33]
port 513 nsew
rlabel metal3 s 0 70456 480 70576 6 gpio_vtrip_sel[34]
port 514 nsew
rlabel metal3 s 0 50872 480 50992 6 gpio_vtrip_sel[35]
port 515 nsew
rlabel metal3 s 0 31288 480 31408 6 gpio_vtrip_sel[36]
port 516 nsew
rlabel metal3 s 0 11704 480 11824 6 gpio_vtrip_sel[37]
port 517 nsew
rlabel metal2 s 37738 0 37794 480 6 gpio_vtrip_sel[38]
port 518 nsew
rlabel metal2 s 87418 0 87474 480 6 gpio_vtrip_sel[39]
port 519 nsew
rlabel metal3 s 439520 76712 440000 76832 6 gpio_vtrip_sel[3]
port 520 nsew
rlabel metal2 s 137098 0 137154 480 6 gpio_vtrip_sel[40]
port 521 nsew
rlabel metal2 s 186778 0 186834 480 6 gpio_vtrip_sel[41]
port 522 nsew
rlabel metal2 s 236458 0 236514 480 6 gpio_vtrip_sel[42]
port 523 nsew
rlabel metal2 s 286138 0 286194 480 6 gpio_vtrip_sel[43]
port 524 nsew
rlabel metal3 s 439520 93032 440000 93152 6 gpio_vtrip_sel[4]
port 525 nsew
rlabel metal3 s 439520 109352 440000 109472 6 gpio_vtrip_sel[5]
port 526 nsew
rlabel metal3 s 439520 125672 440000 125792 6 gpio_vtrip_sel[6]
port 527 nsew
rlabel metal3 s 439520 141992 440000 142112 6 gpio_vtrip_sel[7]
port 528 nsew
rlabel metal3 s 439520 158312 440000 158432 6 gpio_vtrip_sel[8]
port 529 nsew
rlabel metal3 s 439520 174632 440000 174752 6 gpio_vtrip_sel[9]
port 530 nsew
rlabel metal2 s 306838 0 306894 480 6 mask_rev[0]
port 531 nsew
rlabel metal2 s 348238 0 348294 480 6 mask_rev[10]
port 532 nsew
rlabel metal2 s 352378 0 352434 480 6 mask_rev[11]
port 533 nsew
rlabel metal2 s 356518 0 356574 480 6 mask_rev[12]
port 534 nsew
rlabel metal2 s 360658 0 360714 480 6 mask_rev[13]
port 535 nsew
rlabel metal2 s 364798 0 364854 480 6 mask_rev[14]
port 536 nsew
rlabel metal2 s 368938 0 368994 480 6 mask_rev[15]
port 537 nsew
rlabel metal2 s 373078 0 373134 480 6 mask_rev[16]
port 538 nsew
rlabel metal2 s 377218 0 377274 480 6 mask_rev[17]
port 539 nsew
rlabel metal2 s 381358 0 381414 480 6 mask_rev[18]
port 540 nsew
rlabel metal2 s 385498 0 385554 480 6 mask_rev[19]
port 541 nsew
rlabel metal2 s 310978 0 311034 480 6 mask_rev[1]
port 542 nsew
rlabel metal2 s 389638 0 389694 480 6 mask_rev[20]
port 543 nsew
rlabel metal2 s 393778 0 393834 480 6 mask_rev[21]
port 544 nsew
rlabel metal2 s 397918 0 397974 480 6 mask_rev[22]
port 545 nsew
rlabel metal2 s 402058 0 402114 480 6 mask_rev[23]
port 546 nsew
rlabel metal2 s 406198 0 406254 480 6 mask_rev[24]
port 547 nsew
rlabel metal2 s 410338 0 410394 480 6 mask_rev[25]
port 548 nsew
rlabel metal2 s 414478 0 414534 480 6 mask_rev[26]
port 549 nsew
rlabel metal2 s 418618 0 418674 480 6 mask_rev[27]
port 550 nsew
rlabel metal2 s 422758 0 422814 480 6 mask_rev[28]
port 551 nsew
rlabel metal2 s 426898 0 426954 480 6 mask_rev[29]
port 552 nsew
rlabel metal2 s 315118 0 315174 480 6 mask_rev[2]
port 553 nsew
rlabel metal2 s 431038 0 431094 480 6 mask_rev[30]
port 554 nsew
rlabel metal2 s 435178 0 435234 480 6 mask_rev[31]
port 555 nsew
rlabel metal2 s 319258 0 319314 480 6 mask_rev[3]
port 556 nsew
rlabel metal2 s 323398 0 323454 480 6 mask_rev[4]
port 557 nsew
rlabel metal2 s 327538 0 327594 480 6 mask_rev[5]
port 558 nsew
rlabel metal2 s 331678 0 331734 480 6 mask_rev[6]
port 559 nsew
rlabel metal2 s 335818 0 335874 480 6 mask_rev[7]
port 560 nsew
rlabel metal2 s 339958 0 340014 480 6 mask_rev[8]
port 561 nsew
rlabel metal2 s 344098 0 344154 480 6 mask_rev[9]
port 562 nsew
rlabel metal3 s 0 3544 480 3664 6 por
port 563 nsew
rlabel metal3 s 0 1912 480 2032 6 porb
port 564 nsew
rlabel metal2 s 4618 0 4674 480 6 resetb
port 565 nsew
<< properties >>
string FIXED_BBOX 0 0 440000 280000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 182469824
string GDS_FILE /home/karim/work/caravel_openframe_project/openlane/picosoc/runs/picosoc-pll-antenna/results/signoff/picosoc.magic.gds
string GDS_START 17745992
<< end >>

