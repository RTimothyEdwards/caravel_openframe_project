magic
tech sky130A
magscale 1 2
timestamp 1691505922
<< obsli1 >>
rect 1104 2159 438840 297585
<< obsm1 >>
rect 14 1844 439194 298104
<< metal2 >>
rect 3330 299520 3386 300000
rect 7378 299520 7434 300000
rect 11426 299520 11482 300000
rect 15474 299520 15530 300000
rect 19522 299520 19578 300000
rect 23570 299520 23626 300000
rect 27618 299520 27674 300000
rect 31666 299520 31722 300000
rect 35714 299520 35770 300000
rect 39762 299520 39818 300000
rect 43810 299520 43866 300000
rect 47858 299520 47914 300000
rect 51906 299520 51962 300000
rect 55954 299520 56010 300000
rect 60002 299520 60058 300000
rect 64050 299520 64106 300000
rect 68098 299520 68154 300000
rect 72146 299520 72202 300000
rect 76194 299520 76250 300000
rect 80242 299520 80298 300000
rect 84290 299520 84346 300000
rect 88338 299520 88394 300000
rect 92386 299520 92442 300000
rect 96434 299520 96490 300000
rect 100482 299520 100538 300000
rect 104530 299520 104586 300000
rect 108578 299520 108634 300000
rect 112626 299520 112682 300000
rect 116674 299520 116730 300000
rect 120722 299520 120778 300000
rect 124770 299520 124826 300000
rect 128818 299520 128874 300000
rect 132866 299520 132922 300000
rect 136914 299520 136970 300000
rect 140962 299520 141018 300000
rect 145010 299520 145066 300000
rect 149058 299520 149114 300000
rect 153106 299520 153162 300000
rect 157154 299520 157210 300000
rect 161202 299520 161258 300000
rect 165250 299520 165306 300000
rect 169298 299520 169354 300000
rect 173346 299520 173402 300000
rect 177394 299520 177450 300000
rect 181442 299520 181498 300000
rect 185490 299520 185546 300000
rect 189538 299520 189594 300000
rect 193586 299520 193642 300000
rect 197634 299520 197690 300000
rect 201682 299520 201738 300000
rect 205730 299520 205786 300000
rect 209778 299520 209834 300000
rect 213826 299520 213882 300000
rect 217874 299520 217930 300000
rect 221922 299520 221978 300000
rect 225970 299520 226026 300000
rect 230018 299520 230074 300000
rect 234066 299520 234122 300000
rect 238114 299520 238170 300000
rect 242162 299520 242218 300000
rect 246210 299520 246266 300000
rect 250258 299520 250314 300000
rect 254306 299520 254362 300000
rect 258354 299520 258410 300000
rect 262402 299520 262458 300000
rect 266450 299520 266506 300000
rect 270498 299520 270554 300000
rect 274546 299520 274602 300000
rect 278594 299520 278650 300000
rect 282642 299520 282698 300000
rect 286690 299520 286746 300000
rect 290738 299520 290794 300000
rect 294786 299520 294842 300000
rect 298834 299520 298890 300000
rect 302882 299520 302938 300000
rect 306930 299520 306986 300000
rect 310978 299520 311034 300000
rect 315026 299520 315082 300000
rect 319074 299520 319130 300000
rect 323122 299520 323178 300000
rect 327170 299520 327226 300000
rect 331218 299520 331274 300000
rect 335266 299520 335322 300000
rect 339314 299520 339370 300000
rect 343362 299520 343418 300000
rect 347410 299520 347466 300000
rect 351458 299520 351514 300000
rect 355506 299520 355562 300000
rect 359554 299520 359610 300000
rect 363602 299520 363658 300000
rect 367650 299520 367706 300000
rect 371698 299520 371754 300000
rect 375746 299520 375802 300000
rect 379794 299520 379850 300000
rect 383842 299520 383898 300000
rect 387890 299520 387946 300000
rect 391938 299520 391994 300000
rect 395986 299520 396042 300000
rect 400034 299520 400090 300000
rect 404082 299520 404138 300000
rect 408130 299520 408186 300000
rect 412178 299520 412234 300000
rect 416226 299520 416282 300000
rect 420274 299520 420330 300000
rect 424322 299520 424378 300000
rect 428370 299520 428426 300000
rect 432418 299520 432474 300000
rect 436466 299520 436522 300000
rect 4618 0 4674 480
rect 8758 0 8814 480
rect 12898 0 12954 480
rect 17038 0 17094 480
rect 21178 0 21234 480
rect 25318 0 25374 480
rect 29458 0 29514 480
rect 33598 0 33654 480
rect 37738 0 37794 480
rect 41878 0 41934 480
rect 46018 0 46074 480
rect 50158 0 50214 480
rect 54298 0 54354 480
rect 58438 0 58494 480
rect 62578 0 62634 480
rect 66718 0 66774 480
rect 70858 0 70914 480
rect 74998 0 75054 480
rect 79138 0 79194 480
rect 83278 0 83334 480
rect 87418 0 87474 480
rect 91558 0 91614 480
rect 95698 0 95754 480
rect 99838 0 99894 480
rect 103978 0 104034 480
rect 108118 0 108174 480
rect 112258 0 112314 480
rect 116398 0 116454 480
rect 120538 0 120594 480
rect 124678 0 124734 480
rect 128818 0 128874 480
rect 132958 0 133014 480
rect 137098 0 137154 480
rect 141238 0 141294 480
rect 145378 0 145434 480
rect 149518 0 149574 480
rect 153658 0 153714 480
rect 157798 0 157854 480
rect 161938 0 161994 480
rect 166078 0 166134 480
rect 170218 0 170274 480
rect 174358 0 174414 480
rect 178498 0 178554 480
rect 182638 0 182694 480
rect 186778 0 186834 480
rect 190918 0 190974 480
rect 195058 0 195114 480
rect 199198 0 199254 480
rect 203338 0 203394 480
rect 207478 0 207534 480
rect 211618 0 211674 480
rect 215758 0 215814 480
rect 219898 0 219954 480
rect 224038 0 224094 480
rect 228178 0 228234 480
rect 232318 0 232374 480
rect 236458 0 236514 480
rect 240598 0 240654 480
rect 244738 0 244794 480
rect 248878 0 248934 480
rect 253018 0 253074 480
rect 257158 0 257214 480
rect 261298 0 261354 480
rect 265438 0 265494 480
rect 269578 0 269634 480
rect 273718 0 273774 480
rect 277858 0 277914 480
rect 281998 0 282054 480
rect 286138 0 286194 480
rect 290278 0 290334 480
rect 294418 0 294474 480
rect 298558 0 298614 480
rect 302698 0 302754 480
rect 306838 0 306894 480
rect 310978 0 311034 480
rect 315118 0 315174 480
rect 319258 0 319314 480
rect 323398 0 323454 480
rect 327538 0 327594 480
rect 331678 0 331734 480
rect 335818 0 335874 480
rect 339958 0 340014 480
rect 344098 0 344154 480
rect 348238 0 348294 480
rect 352378 0 352434 480
rect 356518 0 356574 480
rect 360658 0 360714 480
rect 364798 0 364854 480
rect 368938 0 368994 480
rect 373078 0 373134 480
rect 377218 0 377274 480
rect 381358 0 381414 480
rect 385498 0 385554 480
rect 389638 0 389694 480
rect 393778 0 393834 480
rect 397918 0 397974 480
rect 402058 0 402114 480
rect 406198 0 406254 480
rect 410338 0 410394 480
rect 414478 0 414534 480
rect 418618 0 418674 480
rect 422758 0 422814 480
rect 426898 0 426954 480
rect 431038 0 431094 480
rect 435178 0 435234 480
<< obsm2 >>
rect 18 299464 3274 299554
rect 3442 299464 7322 299554
rect 7490 299464 11370 299554
rect 11538 299464 15418 299554
rect 15586 299464 19466 299554
rect 19634 299464 23514 299554
rect 23682 299464 27562 299554
rect 27730 299464 31610 299554
rect 31778 299464 35658 299554
rect 35826 299464 39706 299554
rect 39874 299464 43754 299554
rect 43922 299464 47802 299554
rect 47970 299464 51850 299554
rect 52018 299464 55898 299554
rect 56066 299464 59946 299554
rect 60114 299464 63994 299554
rect 64162 299464 68042 299554
rect 68210 299464 72090 299554
rect 72258 299464 76138 299554
rect 76306 299464 80186 299554
rect 80354 299464 84234 299554
rect 84402 299464 88282 299554
rect 88450 299464 92330 299554
rect 92498 299464 96378 299554
rect 96546 299464 100426 299554
rect 100594 299464 104474 299554
rect 104642 299464 108522 299554
rect 108690 299464 112570 299554
rect 112738 299464 116618 299554
rect 116786 299464 120666 299554
rect 120834 299464 124714 299554
rect 124882 299464 128762 299554
rect 128930 299464 132810 299554
rect 132978 299464 136858 299554
rect 137026 299464 140906 299554
rect 141074 299464 144954 299554
rect 145122 299464 149002 299554
rect 149170 299464 153050 299554
rect 153218 299464 157098 299554
rect 157266 299464 161146 299554
rect 161314 299464 165194 299554
rect 165362 299464 169242 299554
rect 169410 299464 173290 299554
rect 173458 299464 177338 299554
rect 177506 299464 181386 299554
rect 181554 299464 185434 299554
rect 185602 299464 189482 299554
rect 189650 299464 193530 299554
rect 193698 299464 197578 299554
rect 197746 299464 201626 299554
rect 201794 299464 205674 299554
rect 205842 299464 209722 299554
rect 209890 299464 213770 299554
rect 213938 299464 217818 299554
rect 217986 299464 221866 299554
rect 222034 299464 225914 299554
rect 226082 299464 229962 299554
rect 230130 299464 234010 299554
rect 234178 299464 238058 299554
rect 238226 299464 242106 299554
rect 242274 299464 246154 299554
rect 246322 299464 250202 299554
rect 250370 299464 254250 299554
rect 254418 299464 258298 299554
rect 258466 299464 262346 299554
rect 262514 299464 266394 299554
rect 266562 299464 270442 299554
rect 270610 299464 274490 299554
rect 274658 299464 278538 299554
rect 278706 299464 282586 299554
rect 282754 299464 286634 299554
rect 286802 299464 290682 299554
rect 290850 299464 294730 299554
rect 294898 299464 298778 299554
rect 298946 299464 302826 299554
rect 302994 299464 306874 299554
rect 307042 299464 310922 299554
rect 311090 299464 314970 299554
rect 315138 299464 319018 299554
rect 319186 299464 323066 299554
rect 323234 299464 327114 299554
rect 327282 299464 331162 299554
rect 331330 299464 335210 299554
rect 335378 299464 339258 299554
rect 339426 299464 343306 299554
rect 343474 299464 347354 299554
rect 347522 299464 351402 299554
rect 351570 299464 355450 299554
rect 355618 299464 359498 299554
rect 359666 299464 363546 299554
rect 363714 299464 367594 299554
rect 367762 299464 371642 299554
rect 371810 299464 375690 299554
rect 375858 299464 379738 299554
rect 379906 299464 383786 299554
rect 383954 299464 387834 299554
rect 388002 299464 391882 299554
rect 392050 299464 395930 299554
rect 396098 299464 399978 299554
rect 400146 299464 404026 299554
rect 404194 299464 408074 299554
rect 408242 299464 412122 299554
rect 412290 299464 416170 299554
rect 416338 299464 420218 299554
rect 420386 299464 424266 299554
rect 424434 299464 428314 299554
rect 428482 299464 432362 299554
rect 432530 299464 436410 299554
rect 436578 299464 439190 299554
rect 18 536 439190 299464
rect 18 326 4562 536
rect 4730 326 8702 536
rect 8870 326 12842 536
rect 13010 326 16982 536
rect 17150 326 21122 536
rect 21290 326 25262 536
rect 25430 326 29402 536
rect 29570 326 33542 536
rect 33710 326 37682 536
rect 37850 326 41822 536
rect 41990 326 45962 536
rect 46130 326 50102 536
rect 50270 326 54242 536
rect 54410 326 58382 536
rect 58550 326 62522 536
rect 62690 326 66662 536
rect 66830 326 70802 536
rect 70970 326 74942 536
rect 75110 326 79082 536
rect 79250 326 83222 536
rect 83390 326 87362 536
rect 87530 326 91502 536
rect 91670 326 95642 536
rect 95810 326 99782 536
rect 99950 326 103922 536
rect 104090 326 108062 536
rect 108230 326 112202 536
rect 112370 326 116342 536
rect 116510 326 120482 536
rect 120650 326 124622 536
rect 124790 326 128762 536
rect 128930 326 132902 536
rect 133070 326 137042 536
rect 137210 326 141182 536
rect 141350 326 145322 536
rect 145490 326 149462 536
rect 149630 326 153602 536
rect 153770 326 157742 536
rect 157910 326 161882 536
rect 162050 326 166022 536
rect 166190 326 170162 536
rect 170330 326 174302 536
rect 174470 326 178442 536
rect 178610 326 182582 536
rect 182750 326 186722 536
rect 186890 326 190862 536
rect 191030 326 195002 536
rect 195170 326 199142 536
rect 199310 326 203282 536
rect 203450 326 207422 536
rect 207590 326 211562 536
rect 211730 326 215702 536
rect 215870 326 219842 536
rect 220010 326 223982 536
rect 224150 326 228122 536
rect 228290 326 232262 536
rect 232430 326 236402 536
rect 236570 326 240542 536
rect 240710 326 244682 536
rect 244850 326 248822 536
rect 248990 326 252962 536
rect 253130 326 257102 536
rect 257270 326 261242 536
rect 261410 326 265382 536
rect 265550 326 269522 536
rect 269690 326 273662 536
rect 273830 326 277802 536
rect 277970 326 281942 536
rect 282110 326 286082 536
rect 286250 326 290222 536
rect 290390 326 294362 536
rect 294530 326 298502 536
rect 298670 326 302642 536
rect 302810 326 306782 536
rect 306950 326 310922 536
rect 311090 326 315062 536
rect 315230 326 319202 536
rect 319370 326 323342 536
rect 323510 326 327482 536
rect 327650 326 331622 536
rect 331790 326 335762 536
rect 335930 326 339902 536
rect 340070 326 344042 536
rect 344210 326 348182 536
rect 348350 326 352322 536
rect 352490 326 356462 536
rect 356630 326 360602 536
rect 360770 326 364742 536
rect 364910 326 368882 536
rect 369050 326 373022 536
rect 373190 326 377162 536
rect 377330 326 381302 536
rect 381470 326 385442 536
rect 385610 326 389582 536
rect 389750 326 393722 536
rect 393890 326 397862 536
rect 398030 326 402002 536
rect 402170 326 406142 536
rect 406310 326 410282 536
rect 410450 326 414422 536
rect 414590 326 418562 536
rect 418730 326 422702 536
rect 422870 326 426842 536
rect 427010 326 430982 536
rect 431150 326 435122 536
rect 435290 326 439190 536
<< metal3 >>
rect 439520 295944 440000 296064
rect 439520 294312 440000 294432
rect 439520 292680 440000 292800
rect 439520 291048 440000 291168
rect 439520 289416 440000 289536
rect 0 287784 480 287904
rect 439520 287784 440000 287904
rect 0 286152 480 286272
rect 439520 286152 440000 286272
rect 0 284520 480 284640
rect 439520 284520 440000 284640
rect 0 282888 480 283008
rect 439520 282888 440000 283008
rect 0 281256 480 281376
rect 439520 281256 440000 281376
rect 0 279624 480 279744
rect 439520 279624 440000 279744
rect 0 277992 480 278112
rect 439520 277992 440000 278112
rect 0 276360 480 276480
rect 439520 276360 440000 276480
rect 0 274728 480 274848
rect 439520 274728 440000 274848
rect 0 273096 480 273216
rect 439520 273096 440000 273216
rect 0 271464 480 271584
rect 439520 271464 440000 271584
rect 0 269832 480 269952
rect 439520 269832 440000 269952
rect 0 268200 480 268320
rect 439520 268200 440000 268320
rect 0 266568 480 266688
rect 439520 266568 440000 266688
rect 0 264936 480 265056
rect 439520 264936 440000 265056
rect 0 263304 480 263424
rect 439520 263304 440000 263424
rect 0 261672 480 261792
rect 439520 261672 440000 261792
rect 0 260040 480 260160
rect 439520 260040 440000 260160
rect 0 258408 480 258528
rect 439520 258408 440000 258528
rect 0 256776 480 256896
rect 439520 256776 440000 256896
rect 0 255144 480 255264
rect 439520 255144 440000 255264
rect 0 253512 480 253632
rect 439520 253512 440000 253632
rect 0 251880 480 252000
rect 439520 251880 440000 252000
rect 0 250248 480 250368
rect 439520 250248 440000 250368
rect 0 248616 480 248736
rect 439520 248616 440000 248736
rect 0 246984 480 247104
rect 439520 246984 440000 247104
rect 0 245352 480 245472
rect 439520 245352 440000 245472
rect 0 243720 480 243840
rect 439520 243720 440000 243840
rect 0 242088 480 242208
rect 439520 242088 440000 242208
rect 0 240456 480 240576
rect 439520 240456 440000 240576
rect 0 238824 480 238944
rect 439520 238824 440000 238944
rect 0 237192 480 237312
rect 439520 237192 440000 237312
rect 0 235560 480 235680
rect 439520 235560 440000 235680
rect 0 233928 480 234048
rect 439520 233928 440000 234048
rect 0 232296 480 232416
rect 439520 232296 440000 232416
rect 0 230664 480 230784
rect 439520 230664 440000 230784
rect 0 229032 480 229152
rect 439520 229032 440000 229152
rect 0 227400 480 227520
rect 439520 227400 440000 227520
rect 0 225768 480 225888
rect 439520 225768 440000 225888
rect 0 224136 480 224256
rect 439520 224136 440000 224256
rect 0 222504 480 222624
rect 439520 222504 440000 222624
rect 0 220872 480 220992
rect 439520 220872 440000 220992
rect 0 219240 480 219360
rect 439520 219240 440000 219360
rect 0 217608 480 217728
rect 439520 217608 440000 217728
rect 0 215976 480 216096
rect 439520 215976 440000 216096
rect 0 214344 480 214464
rect 439520 214344 440000 214464
rect 0 212712 480 212832
rect 439520 212712 440000 212832
rect 0 211080 480 211200
rect 439520 211080 440000 211200
rect 0 209448 480 209568
rect 439520 209448 440000 209568
rect 0 207816 480 207936
rect 439520 207816 440000 207936
rect 0 206184 480 206304
rect 439520 206184 440000 206304
rect 0 204552 480 204672
rect 439520 204552 440000 204672
rect 0 202920 480 203040
rect 439520 202920 440000 203040
rect 0 201288 480 201408
rect 439520 201288 440000 201408
rect 0 199656 480 199776
rect 439520 199656 440000 199776
rect 0 198024 480 198144
rect 439520 198024 440000 198144
rect 0 196392 480 196512
rect 439520 196392 440000 196512
rect 0 194760 480 194880
rect 439520 194760 440000 194880
rect 0 193128 480 193248
rect 439520 193128 440000 193248
rect 0 191496 480 191616
rect 439520 191496 440000 191616
rect 0 189864 480 189984
rect 439520 189864 440000 189984
rect 0 188232 480 188352
rect 439520 188232 440000 188352
rect 0 186600 480 186720
rect 439520 186600 440000 186720
rect 0 184968 480 185088
rect 439520 184968 440000 185088
rect 0 183336 480 183456
rect 439520 183336 440000 183456
rect 0 181704 480 181824
rect 439520 181704 440000 181824
rect 0 180072 480 180192
rect 439520 180072 440000 180192
rect 0 178440 480 178560
rect 439520 178440 440000 178560
rect 0 176808 480 176928
rect 439520 176808 440000 176928
rect 0 175176 480 175296
rect 439520 175176 440000 175296
rect 0 173544 480 173664
rect 439520 173544 440000 173664
rect 0 171912 480 172032
rect 439520 171912 440000 172032
rect 0 170280 480 170400
rect 439520 170280 440000 170400
rect 0 168648 480 168768
rect 439520 168648 440000 168768
rect 0 167016 480 167136
rect 439520 167016 440000 167136
rect 0 165384 480 165504
rect 439520 165384 440000 165504
rect 0 163752 480 163872
rect 439520 163752 440000 163872
rect 0 162120 480 162240
rect 439520 162120 440000 162240
rect 0 160488 480 160608
rect 439520 160488 440000 160608
rect 0 158856 480 158976
rect 439520 158856 440000 158976
rect 0 157224 480 157344
rect 439520 157224 440000 157344
rect 0 155592 480 155712
rect 439520 155592 440000 155712
rect 0 153960 480 154080
rect 439520 153960 440000 154080
rect 0 152328 480 152448
rect 439520 152328 440000 152448
rect 0 150696 480 150816
rect 439520 150696 440000 150816
rect 0 149064 480 149184
rect 439520 149064 440000 149184
rect 0 147432 480 147552
rect 439520 147432 440000 147552
rect 0 145800 480 145920
rect 439520 145800 440000 145920
rect 0 144168 480 144288
rect 439520 144168 440000 144288
rect 0 142536 480 142656
rect 439520 142536 440000 142656
rect 0 140904 480 141024
rect 439520 140904 440000 141024
rect 0 139272 480 139392
rect 439520 139272 440000 139392
rect 0 137640 480 137760
rect 439520 137640 440000 137760
rect 0 136008 480 136128
rect 439520 136008 440000 136128
rect 0 134376 480 134496
rect 439520 134376 440000 134496
rect 0 132744 480 132864
rect 439520 132744 440000 132864
rect 0 131112 480 131232
rect 439520 131112 440000 131232
rect 0 129480 480 129600
rect 439520 129480 440000 129600
rect 0 127848 480 127968
rect 439520 127848 440000 127968
rect 0 126216 480 126336
rect 439520 126216 440000 126336
rect 0 124584 480 124704
rect 439520 124584 440000 124704
rect 0 122952 480 123072
rect 439520 122952 440000 123072
rect 0 121320 480 121440
rect 439520 121320 440000 121440
rect 0 119688 480 119808
rect 439520 119688 440000 119808
rect 0 118056 480 118176
rect 439520 118056 440000 118176
rect 0 116424 480 116544
rect 439520 116424 440000 116544
rect 0 114792 480 114912
rect 439520 114792 440000 114912
rect 0 113160 480 113280
rect 439520 113160 440000 113280
rect 0 111528 480 111648
rect 439520 111528 440000 111648
rect 0 109896 480 110016
rect 439520 109896 440000 110016
rect 0 108264 480 108384
rect 439520 108264 440000 108384
rect 0 106632 480 106752
rect 439520 106632 440000 106752
rect 0 105000 480 105120
rect 439520 105000 440000 105120
rect 0 103368 480 103488
rect 439520 103368 440000 103488
rect 0 101736 480 101856
rect 439520 101736 440000 101856
rect 0 100104 480 100224
rect 439520 100104 440000 100224
rect 0 98472 480 98592
rect 439520 98472 440000 98592
rect 0 96840 480 96960
rect 439520 96840 440000 96960
rect 0 95208 480 95328
rect 439520 95208 440000 95328
rect 0 93576 480 93696
rect 439520 93576 440000 93696
rect 0 91944 480 92064
rect 439520 91944 440000 92064
rect 0 90312 480 90432
rect 439520 90312 440000 90432
rect 0 88680 480 88800
rect 439520 88680 440000 88800
rect 0 87048 480 87168
rect 439520 87048 440000 87168
rect 0 85416 480 85536
rect 439520 85416 440000 85536
rect 0 83784 480 83904
rect 439520 83784 440000 83904
rect 0 82152 480 82272
rect 439520 82152 440000 82272
rect 0 80520 480 80640
rect 439520 80520 440000 80640
rect 0 78888 480 79008
rect 439520 78888 440000 79008
rect 0 77256 480 77376
rect 439520 77256 440000 77376
rect 0 75624 480 75744
rect 439520 75624 440000 75744
rect 0 73992 480 74112
rect 439520 73992 440000 74112
rect 0 72360 480 72480
rect 439520 72360 440000 72480
rect 0 70728 480 70848
rect 439520 70728 440000 70848
rect 0 69096 480 69216
rect 439520 69096 440000 69216
rect 0 67464 480 67584
rect 439520 67464 440000 67584
rect 0 65832 480 65952
rect 439520 65832 440000 65952
rect 0 64200 480 64320
rect 439520 64200 440000 64320
rect 0 62568 480 62688
rect 439520 62568 440000 62688
rect 0 60936 480 61056
rect 439520 60936 440000 61056
rect 0 59304 480 59424
rect 439520 59304 440000 59424
rect 0 57672 480 57792
rect 439520 57672 440000 57792
rect 0 56040 480 56160
rect 439520 56040 440000 56160
rect 0 54408 480 54528
rect 439520 54408 440000 54528
rect 0 52776 480 52896
rect 439520 52776 440000 52896
rect 0 51144 480 51264
rect 439520 51144 440000 51264
rect 0 49512 480 49632
rect 439520 49512 440000 49632
rect 0 47880 480 48000
rect 439520 47880 440000 48000
rect 0 46248 480 46368
rect 439520 46248 440000 46368
rect 0 44616 480 44736
rect 439520 44616 440000 44736
rect 0 42984 480 43104
rect 439520 42984 440000 43104
rect 0 41352 480 41472
rect 439520 41352 440000 41472
rect 0 39720 480 39840
rect 439520 39720 440000 39840
rect 0 38088 480 38208
rect 439520 38088 440000 38208
rect 0 36456 480 36576
rect 439520 36456 440000 36576
rect 0 34824 480 34944
rect 439520 34824 440000 34944
rect 0 33192 480 33312
rect 439520 33192 440000 33312
rect 0 31560 480 31680
rect 439520 31560 440000 31680
rect 0 29928 480 30048
rect 439520 29928 440000 30048
rect 0 28296 480 28416
rect 439520 28296 440000 28416
rect 0 26664 480 26784
rect 439520 26664 440000 26784
rect 0 25032 480 25152
rect 439520 25032 440000 25152
rect 0 23400 480 23520
rect 439520 23400 440000 23520
rect 0 21768 480 21888
rect 439520 21768 440000 21888
rect 0 20136 480 20256
rect 439520 20136 440000 20256
rect 0 18504 480 18624
rect 439520 18504 440000 18624
rect 0 16872 480 16992
rect 439520 16872 440000 16992
rect 0 15240 480 15360
rect 439520 15240 440000 15360
rect 0 13608 480 13728
rect 439520 13608 440000 13728
rect 0 11976 480 12096
rect 439520 11976 440000 12096
rect 439520 10344 440000 10464
rect 439520 8712 440000 8832
rect 439520 7080 440000 7200
rect 439520 5448 440000 5568
rect 439520 3816 440000 3936
<< obsm3 >>
rect 480 296144 439520 297601
rect 480 295864 439440 296144
rect 480 294512 439520 295864
rect 480 294232 439440 294512
rect 480 292880 439520 294232
rect 480 292600 439440 292880
rect 480 291248 439520 292600
rect 480 290968 439440 291248
rect 480 289616 439520 290968
rect 480 289336 439440 289616
rect 480 287984 439520 289336
rect 560 287704 439440 287984
rect 480 286352 439520 287704
rect 560 286072 439440 286352
rect 480 284720 439520 286072
rect 560 284440 439440 284720
rect 480 283088 439520 284440
rect 560 282808 439440 283088
rect 480 281456 439520 282808
rect 560 281176 439440 281456
rect 480 279824 439520 281176
rect 560 279544 439440 279824
rect 480 278192 439520 279544
rect 560 277912 439440 278192
rect 480 276560 439520 277912
rect 560 276280 439440 276560
rect 480 274928 439520 276280
rect 560 274648 439440 274928
rect 480 273296 439520 274648
rect 560 273016 439440 273296
rect 480 271664 439520 273016
rect 560 271384 439440 271664
rect 480 270032 439520 271384
rect 560 269752 439440 270032
rect 480 268400 439520 269752
rect 560 268120 439440 268400
rect 480 266768 439520 268120
rect 560 266488 439440 266768
rect 480 265136 439520 266488
rect 560 264856 439440 265136
rect 480 263504 439520 264856
rect 560 263224 439440 263504
rect 480 261872 439520 263224
rect 560 261592 439440 261872
rect 480 260240 439520 261592
rect 560 259960 439440 260240
rect 480 258608 439520 259960
rect 560 258328 439440 258608
rect 480 256976 439520 258328
rect 560 256696 439440 256976
rect 480 255344 439520 256696
rect 560 255064 439440 255344
rect 480 253712 439520 255064
rect 560 253432 439440 253712
rect 480 252080 439520 253432
rect 560 251800 439440 252080
rect 480 250448 439520 251800
rect 560 250168 439440 250448
rect 480 248816 439520 250168
rect 560 248536 439440 248816
rect 480 247184 439520 248536
rect 560 246904 439440 247184
rect 480 245552 439520 246904
rect 560 245272 439440 245552
rect 480 243920 439520 245272
rect 560 243640 439440 243920
rect 480 242288 439520 243640
rect 560 242008 439440 242288
rect 480 240656 439520 242008
rect 560 240376 439440 240656
rect 480 239024 439520 240376
rect 560 238744 439440 239024
rect 480 237392 439520 238744
rect 560 237112 439440 237392
rect 480 235760 439520 237112
rect 560 235480 439440 235760
rect 480 234128 439520 235480
rect 560 233848 439440 234128
rect 480 232496 439520 233848
rect 560 232216 439440 232496
rect 480 230864 439520 232216
rect 560 230584 439440 230864
rect 480 229232 439520 230584
rect 560 228952 439440 229232
rect 480 227600 439520 228952
rect 560 227320 439440 227600
rect 480 225968 439520 227320
rect 560 225688 439440 225968
rect 480 224336 439520 225688
rect 560 224056 439440 224336
rect 480 222704 439520 224056
rect 560 222424 439440 222704
rect 480 221072 439520 222424
rect 560 220792 439440 221072
rect 480 219440 439520 220792
rect 560 219160 439440 219440
rect 480 217808 439520 219160
rect 560 217528 439440 217808
rect 480 216176 439520 217528
rect 560 215896 439440 216176
rect 480 214544 439520 215896
rect 560 214264 439440 214544
rect 480 212912 439520 214264
rect 560 212632 439440 212912
rect 480 211280 439520 212632
rect 560 211000 439440 211280
rect 480 209648 439520 211000
rect 560 209368 439440 209648
rect 480 208016 439520 209368
rect 560 207736 439440 208016
rect 480 206384 439520 207736
rect 560 206104 439440 206384
rect 480 204752 439520 206104
rect 560 204472 439440 204752
rect 480 203120 439520 204472
rect 560 202840 439440 203120
rect 480 201488 439520 202840
rect 560 201208 439440 201488
rect 480 199856 439520 201208
rect 560 199576 439440 199856
rect 480 198224 439520 199576
rect 560 197944 439440 198224
rect 480 196592 439520 197944
rect 560 196312 439440 196592
rect 480 194960 439520 196312
rect 560 194680 439440 194960
rect 480 193328 439520 194680
rect 560 193048 439440 193328
rect 480 191696 439520 193048
rect 560 191416 439440 191696
rect 480 190064 439520 191416
rect 560 189784 439440 190064
rect 480 188432 439520 189784
rect 560 188152 439440 188432
rect 480 186800 439520 188152
rect 560 186520 439440 186800
rect 480 185168 439520 186520
rect 560 184888 439440 185168
rect 480 183536 439520 184888
rect 560 183256 439440 183536
rect 480 181904 439520 183256
rect 560 181624 439440 181904
rect 480 180272 439520 181624
rect 560 179992 439440 180272
rect 480 178640 439520 179992
rect 560 178360 439440 178640
rect 480 177008 439520 178360
rect 560 176728 439440 177008
rect 480 175376 439520 176728
rect 560 175096 439440 175376
rect 480 173744 439520 175096
rect 560 173464 439440 173744
rect 480 172112 439520 173464
rect 560 171832 439440 172112
rect 480 170480 439520 171832
rect 560 170200 439440 170480
rect 480 168848 439520 170200
rect 560 168568 439440 168848
rect 480 167216 439520 168568
rect 560 166936 439440 167216
rect 480 165584 439520 166936
rect 560 165304 439440 165584
rect 480 163952 439520 165304
rect 560 163672 439440 163952
rect 480 162320 439520 163672
rect 560 162040 439440 162320
rect 480 160688 439520 162040
rect 560 160408 439440 160688
rect 480 159056 439520 160408
rect 560 158776 439440 159056
rect 480 157424 439520 158776
rect 560 157144 439440 157424
rect 480 155792 439520 157144
rect 560 155512 439440 155792
rect 480 154160 439520 155512
rect 560 153880 439440 154160
rect 480 152528 439520 153880
rect 560 152248 439440 152528
rect 480 150896 439520 152248
rect 560 150616 439440 150896
rect 480 149264 439520 150616
rect 560 148984 439440 149264
rect 480 147632 439520 148984
rect 560 147352 439440 147632
rect 480 146000 439520 147352
rect 560 145720 439440 146000
rect 480 144368 439520 145720
rect 560 144088 439440 144368
rect 480 142736 439520 144088
rect 560 142456 439440 142736
rect 480 141104 439520 142456
rect 560 140824 439440 141104
rect 480 139472 439520 140824
rect 560 139192 439440 139472
rect 480 137840 439520 139192
rect 560 137560 439440 137840
rect 480 136208 439520 137560
rect 560 135928 439440 136208
rect 480 134576 439520 135928
rect 560 134296 439440 134576
rect 480 132944 439520 134296
rect 560 132664 439440 132944
rect 480 131312 439520 132664
rect 560 131032 439440 131312
rect 480 129680 439520 131032
rect 560 129400 439440 129680
rect 480 128048 439520 129400
rect 560 127768 439440 128048
rect 480 126416 439520 127768
rect 560 126136 439440 126416
rect 480 124784 439520 126136
rect 560 124504 439440 124784
rect 480 123152 439520 124504
rect 560 122872 439440 123152
rect 480 121520 439520 122872
rect 560 121240 439440 121520
rect 480 119888 439520 121240
rect 560 119608 439440 119888
rect 480 118256 439520 119608
rect 560 117976 439440 118256
rect 480 116624 439520 117976
rect 560 116344 439440 116624
rect 480 114992 439520 116344
rect 560 114712 439440 114992
rect 480 113360 439520 114712
rect 560 113080 439440 113360
rect 480 111728 439520 113080
rect 560 111448 439440 111728
rect 480 110096 439520 111448
rect 560 109816 439440 110096
rect 480 108464 439520 109816
rect 560 108184 439440 108464
rect 480 106832 439520 108184
rect 560 106552 439440 106832
rect 480 105200 439520 106552
rect 560 104920 439440 105200
rect 480 103568 439520 104920
rect 560 103288 439440 103568
rect 480 101936 439520 103288
rect 560 101656 439440 101936
rect 480 100304 439520 101656
rect 560 100024 439440 100304
rect 480 98672 439520 100024
rect 560 98392 439440 98672
rect 480 97040 439520 98392
rect 560 96760 439440 97040
rect 480 95408 439520 96760
rect 560 95128 439440 95408
rect 480 93776 439520 95128
rect 560 93496 439440 93776
rect 480 92144 439520 93496
rect 560 91864 439440 92144
rect 480 90512 439520 91864
rect 560 90232 439440 90512
rect 480 88880 439520 90232
rect 560 88600 439440 88880
rect 480 87248 439520 88600
rect 560 86968 439440 87248
rect 480 85616 439520 86968
rect 560 85336 439440 85616
rect 480 83984 439520 85336
rect 560 83704 439440 83984
rect 480 82352 439520 83704
rect 560 82072 439440 82352
rect 480 80720 439520 82072
rect 560 80440 439440 80720
rect 480 79088 439520 80440
rect 560 78808 439440 79088
rect 480 77456 439520 78808
rect 560 77176 439440 77456
rect 480 75824 439520 77176
rect 560 75544 439440 75824
rect 480 74192 439520 75544
rect 560 73912 439440 74192
rect 480 72560 439520 73912
rect 560 72280 439440 72560
rect 480 70928 439520 72280
rect 560 70648 439440 70928
rect 480 69296 439520 70648
rect 560 69016 439440 69296
rect 480 67664 439520 69016
rect 560 67384 439440 67664
rect 480 66032 439520 67384
rect 560 65752 439440 66032
rect 480 64400 439520 65752
rect 560 64120 439440 64400
rect 480 62768 439520 64120
rect 560 62488 439440 62768
rect 480 61136 439520 62488
rect 560 60856 439440 61136
rect 480 59504 439520 60856
rect 560 59224 439440 59504
rect 480 57872 439520 59224
rect 560 57592 439440 57872
rect 480 56240 439520 57592
rect 560 55960 439440 56240
rect 480 54608 439520 55960
rect 560 54328 439440 54608
rect 480 52976 439520 54328
rect 560 52696 439440 52976
rect 480 51344 439520 52696
rect 560 51064 439440 51344
rect 480 49712 439520 51064
rect 560 49432 439440 49712
rect 480 48080 439520 49432
rect 560 47800 439440 48080
rect 480 46448 439520 47800
rect 560 46168 439440 46448
rect 480 44816 439520 46168
rect 560 44536 439440 44816
rect 480 43184 439520 44536
rect 560 42904 439440 43184
rect 480 41552 439520 42904
rect 560 41272 439440 41552
rect 480 39920 439520 41272
rect 560 39640 439440 39920
rect 480 38288 439520 39640
rect 560 38008 439440 38288
rect 480 36656 439520 38008
rect 560 36376 439440 36656
rect 480 35024 439520 36376
rect 560 34744 439440 35024
rect 480 33392 439520 34744
rect 560 33112 439440 33392
rect 480 31760 439520 33112
rect 560 31480 439440 31760
rect 480 30128 439520 31480
rect 560 29848 439440 30128
rect 480 28496 439520 29848
rect 560 28216 439440 28496
rect 480 26864 439520 28216
rect 560 26584 439440 26864
rect 480 25232 439520 26584
rect 560 24952 439440 25232
rect 480 23600 439520 24952
rect 560 23320 439440 23600
rect 480 21968 439520 23320
rect 560 21688 439440 21968
rect 480 20336 439520 21688
rect 560 20056 439440 20336
rect 480 18704 439520 20056
rect 560 18424 439440 18704
rect 480 17072 439520 18424
rect 560 16792 439440 17072
rect 480 15440 439520 16792
rect 560 15160 439440 15440
rect 480 13808 439520 15160
rect 560 13528 439440 13808
rect 480 12176 439520 13528
rect 560 11896 439440 12176
rect 480 10544 439520 11896
rect 480 10264 439440 10544
rect 480 8912 439520 10264
rect 480 8632 439440 8912
rect 480 7280 439520 8632
rect 480 7000 439440 7280
rect 480 5648 439520 7000
rect 480 5368 439440 5648
rect 480 4016 439520 5368
rect 480 3736 439440 4016
rect 480 2143 439520 3736
<< metal4 >>
rect 1794 2128 2414 297616
rect 2814 2128 3434 297616
rect 9794 2128 10414 297616
rect 10814 2128 11434 297616
rect 17794 209324 18414 297616
rect 18814 209324 19434 297616
rect 25794 209324 26414 297616
rect 26814 209324 27434 297616
rect 33794 209324 34414 297616
rect 34814 209324 35434 297616
rect 41794 209324 42414 297616
rect 42814 209324 43434 297616
rect 49794 209324 50414 297616
rect 50814 209448 51434 297616
rect 57794 209392 58414 297616
rect 58814 209324 59434 297616
rect 65794 209392 66414 297616
rect 66814 209324 67434 297616
rect 73794 209324 74414 297616
rect 74814 209324 75434 297616
rect 81794 209324 82414 297616
rect 82814 209324 83434 297616
rect 89794 209324 90414 297616
rect 90814 209448 91434 297616
rect 97794 209324 98414 297616
rect 98814 209324 99434 297616
rect 105794 209392 106414 297616
rect 106814 209324 107434 297616
rect 113794 209324 114414 297616
rect 114814 209324 115434 297616
rect 121794 209324 122414 297616
rect 122814 209448 123434 297616
rect 129794 209324 130414 297616
rect 130814 209324 131434 297616
rect 137794 209392 138414 297616
rect 138814 209324 139434 297616
rect 145794 209324 146414 297616
rect 146814 209324 147434 297616
rect 153794 209324 154414 297616
rect 154814 209324 155434 297616
rect 17794 2128 18414 121984
rect 18814 2128 19434 121984
rect 25794 2128 26414 121984
rect 26814 2128 27434 121984
rect 33794 2128 34414 121984
rect 34814 2128 35434 121984
rect 41794 2128 42414 121860
rect 42814 2128 43434 121904
rect 49794 2128 50414 121860
rect 50814 2128 51434 121904
rect 57794 2128 58414 121860
rect 58814 2128 59434 121904
rect 65794 2128 66414 121860
rect 66814 2128 67434 121904
rect 73794 2128 74414 121860
rect 74814 2128 75434 121984
rect 81794 2128 82414 121984
rect 82814 2128 83434 121904
rect 89794 2128 90414 121984
rect 90814 2128 91434 121904
rect 97794 2128 98414 121860
rect 98814 2128 99434 121984
rect 105794 2128 106414 121860
rect 106814 2128 107434 121984
rect 113794 2128 114414 121984
rect 114814 2128 115434 121984
rect 121794 2128 122414 121984
rect 122814 2128 123434 121904
rect 129794 2128 130414 121984
rect 130814 2128 131434 121984
rect 137794 2128 138414 121984
rect 138814 2128 139434 121984
rect 145794 2128 146414 121984
rect 146814 2128 147434 121984
rect 153794 2128 154414 121984
rect 154814 2128 155434 121984
rect 161794 2128 162414 297616
rect 162814 2128 163434 297616
rect 169794 2128 170414 297616
rect 170814 2128 171434 297616
rect 177794 2128 178414 297616
rect 178814 2128 179434 297616
rect 185794 2128 186414 297616
rect 186814 2128 187434 297616
rect 193794 2128 194414 297616
rect 194814 2128 195434 297616
rect 201794 2128 202414 297616
rect 202814 2128 203434 297616
rect 209794 2128 210414 297616
rect 210814 2128 211434 297616
rect 217794 2128 218414 297616
rect 218814 2128 219434 297616
rect 225794 2128 226414 297616
rect 226814 2128 227434 297616
rect 233794 2128 234414 297616
rect 234814 2128 235434 297616
rect 241794 54788 242414 297616
rect 242814 53073 243434 297616
rect 249794 54788 250414 297616
rect 241794 2128 242414 37900
rect 242814 2128 243434 47231
rect 249794 2128 250414 37900
rect 250814 2128 251434 297616
rect 257794 2128 258414 297616
rect 258814 2128 259434 297616
rect 265794 2128 266414 297616
rect 266814 2128 267434 297616
rect 273794 2128 274414 297616
rect 274814 2128 275434 297616
rect 281794 209324 282414 297616
rect 282814 209324 283434 297616
rect 289794 209324 290414 297616
rect 290814 209324 291434 297616
rect 297794 209324 298414 297616
rect 298814 209324 299434 297616
rect 305794 209324 306414 297616
rect 306814 209324 307434 297616
rect 313794 209324 314414 297616
rect 314814 209324 315434 297616
rect 321794 209324 322414 297616
rect 322814 209448 323434 297616
rect 329794 209324 330414 297616
rect 330814 209448 331434 297616
rect 337794 209392 338414 297616
rect 338814 209324 339434 297616
rect 345794 209392 346414 297616
rect 346814 209324 347434 297616
rect 353794 209324 354414 297616
rect 354814 209324 355434 297616
rect 361794 209324 362414 297616
rect 362814 209448 363434 297616
rect 369794 209324 370414 297616
rect 370814 209448 371434 297616
rect 377794 209392 378414 297616
rect 378814 209324 379434 297616
rect 385794 209392 386414 297616
rect 386814 209324 387434 297616
rect 393794 209324 394414 297616
rect 394814 209324 395434 297616
rect 401794 209324 402414 297616
rect 402814 209324 403434 297616
rect 409794 209324 410414 297616
rect 410814 209448 411434 297616
rect 417794 209324 418414 297616
rect 281794 2128 282414 121984
rect 282814 2128 283434 121984
rect 289794 2128 290414 121984
rect 290814 2128 291434 121984
rect 297794 2128 298414 121860
rect 298814 2128 299434 121904
rect 305794 2128 306414 121860
rect 306814 2128 307434 121984
rect 313794 2128 314414 121860
rect 314814 2128 315434 121984
rect 321794 2128 322414 121860
rect 322814 2128 323434 121904
rect 329794 2128 330414 121860
rect 330814 2128 331434 121904
rect 337794 2128 338414 121860
rect 338814 2128 339434 121904
rect 345794 2128 346414 121860
rect 346814 2128 347434 121984
rect 353794 2128 354414 121984
rect 354814 2128 355434 121984
rect 361794 2128 362414 121984
rect 362814 2128 363434 121904
rect 369794 2128 370414 121984
rect 370814 2128 371434 121904
rect 377794 2128 378414 121860
rect 378814 2128 379434 121984
rect 385794 2128 386414 121860
rect 386814 2128 387434 121984
rect 393794 2128 394414 121984
rect 394814 2128 395434 121984
rect 401794 2128 402414 121984
rect 402814 2128 403434 121904
rect 409794 2128 410414 121984
rect 410814 2128 411434 121984
rect 417794 2128 418414 121984
rect 418814 2128 419434 297616
rect 425794 2128 426414 297616
rect 426814 2128 427434 297616
rect 433794 2128 434414 297616
rect 434814 2128 435434 297616
<< obsm4 >>
rect 3739 8195 9714 294677
rect 10494 8195 10734 294677
rect 11514 209244 17714 294677
rect 18494 209244 18734 294677
rect 19514 209244 25714 294677
rect 26494 209244 26734 294677
rect 27514 209244 33714 294677
rect 34494 209244 34734 294677
rect 35514 209244 41714 294677
rect 42494 209244 42734 294677
rect 43514 209244 49714 294677
rect 50494 209368 50734 294677
rect 51514 209368 57714 294677
rect 50494 209312 57714 209368
rect 58494 209312 58734 294677
rect 50494 209244 58734 209312
rect 59514 209312 65714 294677
rect 66494 209312 66734 294677
rect 59514 209244 66734 209312
rect 67514 209244 73714 294677
rect 74494 209244 74734 294677
rect 75514 209244 81714 294677
rect 82494 209244 82734 294677
rect 83514 209244 89714 294677
rect 90494 209368 90734 294677
rect 91514 209368 97714 294677
rect 90494 209244 97714 209368
rect 98494 209244 98734 294677
rect 99514 209312 105714 294677
rect 106494 209312 106734 294677
rect 99514 209244 106734 209312
rect 107514 209244 113714 294677
rect 114494 209244 114734 294677
rect 115514 209244 121714 294677
rect 122494 209368 122734 294677
rect 123514 209368 129714 294677
rect 122494 209244 129714 209368
rect 130494 209244 130734 294677
rect 131514 209312 137714 294677
rect 138494 209312 138734 294677
rect 131514 209244 138734 209312
rect 139514 209244 145714 294677
rect 146494 209244 146734 294677
rect 147514 209244 153714 294677
rect 154494 209244 154734 294677
rect 155514 209244 161714 294677
rect 11514 122064 161714 209244
rect 11514 8195 17714 122064
rect 18494 8195 18734 122064
rect 19514 8195 25714 122064
rect 26494 8195 26734 122064
rect 27514 8195 33714 122064
rect 34494 8195 34734 122064
rect 35514 121984 74734 122064
rect 35514 121940 42734 121984
rect 35514 8195 41714 121940
rect 42494 8195 42734 121940
rect 43514 121940 50734 121984
rect 43514 8195 49714 121940
rect 50494 8195 50734 121940
rect 51514 121940 58734 121984
rect 51514 8195 57714 121940
rect 58494 8195 58734 121940
rect 59514 121940 66734 121984
rect 59514 8195 65714 121940
rect 66494 8195 66734 121940
rect 67514 121940 74734 121984
rect 67514 8195 73714 121940
rect 74494 8195 74734 121940
rect 75514 8195 81714 122064
rect 82494 121984 89714 122064
rect 90494 121984 98734 122064
rect 82494 8195 82734 121984
rect 83514 8195 89714 121984
rect 90494 8195 90734 121984
rect 91514 121940 98734 121984
rect 91514 8195 97714 121940
rect 98494 8195 98734 121940
rect 99514 121940 106734 122064
rect 99514 8195 105714 121940
rect 106494 8195 106734 121940
rect 107514 8195 113714 122064
rect 114494 8195 114734 122064
rect 115514 8195 121714 122064
rect 122494 121984 129714 122064
rect 122494 8195 122734 121984
rect 123514 8195 129714 121984
rect 130494 8195 130734 122064
rect 131514 8195 137714 122064
rect 138494 8195 138734 122064
rect 139514 8195 145714 122064
rect 146494 8195 146734 122064
rect 147514 8195 153714 122064
rect 154494 8195 154734 122064
rect 155514 8195 161714 122064
rect 162494 8195 162734 294677
rect 163514 8195 169714 294677
rect 170494 8195 170734 294677
rect 171514 8195 177714 294677
rect 178494 8195 178734 294677
rect 179514 8195 185714 294677
rect 186494 8195 186734 294677
rect 187514 8195 193714 294677
rect 194494 8195 194734 294677
rect 195514 8195 201714 294677
rect 202494 8195 202734 294677
rect 203514 8195 209714 294677
rect 210494 8195 210734 294677
rect 211514 8195 217714 294677
rect 218494 8195 218734 294677
rect 219514 8195 225714 294677
rect 226494 8195 226734 294677
rect 227514 8195 233714 294677
rect 234494 8195 234734 294677
rect 235514 54708 241714 294677
rect 242494 54708 242734 294677
rect 235514 52993 242734 54708
rect 243514 54708 249714 294677
rect 250494 54708 250734 294677
rect 243514 52993 250734 54708
rect 235514 47311 250734 52993
rect 235514 37980 242734 47311
rect 235514 8195 241714 37980
rect 242494 8195 242734 37980
rect 243514 37980 250734 47311
rect 243514 8195 249714 37980
rect 250494 8195 250734 37980
rect 251514 8195 257714 294677
rect 258494 8195 258734 294677
rect 259514 8195 265714 294677
rect 266494 8195 266734 294677
rect 267514 8195 273714 294677
rect 274494 8195 274734 294677
rect 275514 209244 281714 294677
rect 282494 209244 282734 294677
rect 283514 209244 289714 294677
rect 290494 209244 290734 294677
rect 291514 209244 297714 294677
rect 298494 209244 298734 294677
rect 299514 209244 305714 294677
rect 306494 209244 306734 294677
rect 307514 209244 313714 294677
rect 314494 209244 314734 294677
rect 315514 209244 321714 294677
rect 322494 209368 322734 294677
rect 323514 209368 329714 294677
rect 322494 209244 329714 209368
rect 330494 209368 330734 294677
rect 331514 209368 337714 294677
rect 330494 209312 337714 209368
rect 338494 209312 338734 294677
rect 330494 209244 338734 209312
rect 339514 209312 345714 294677
rect 346494 209312 346734 294677
rect 339514 209244 346734 209312
rect 347514 209244 353714 294677
rect 354494 209244 354734 294677
rect 355514 209244 361714 294677
rect 362494 209368 362734 294677
rect 363514 209368 369714 294677
rect 362494 209244 369714 209368
rect 370494 209368 370734 294677
rect 371514 209368 377714 294677
rect 370494 209312 377714 209368
rect 378494 209312 378734 294677
rect 370494 209244 378734 209312
rect 379514 209312 385714 294677
rect 386494 209312 386734 294677
rect 379514 209244 386734 209312
rect 387514 209244 393714 294677
rect 394494 209244 394734 294677
rect 395514 209244 401714 294677
rect 402494 209244 402734 294677
rect 403514 209244 409714 294677
rect 410494 209368 410734 294677
rect 411514 209368 417714 294677
rect 410494 209244 417714 209368
rect 418494 209244 418734 294677
rect 275514 122064 418734 209244
rect 275514 8195 281714 122064
rect 282494 8195 282734 122064
rect 283514 8195 289714 122064
rect 290494 8195 290734 122064
rect 291514 121984 306734 122064
rect 291514 121940 298734 121984
rect 291514 8195 297714 121940
rect 298494 8195 298734 121940
rect 299514 121940 306734 121984
rect 299514 8195 305714 121940
rect 306494 8195 306734 121940
rect 307514 121940 314734 122064
rect 315514 121984 346734 122064
rect 307514 8195 313714 121940
rect 314494 8195 314734 121940
rect 315514 121940 322734 121984
rect 315514 8195 321714 121940
rect 322494 8195 322734 121940
rect 323514 121940 330734 121984
rect 323514 8195 329714 121940
rect 330494 8195 330734 121940
rect 331514 121940 338734 121984
rect 331514 8195 337714 121940
rect 338494 8195 338734 121940
rect 339514 121940 346734 121984
rect 339514 8195 345714 121940
rect 346494 8195 346734 121940
rect 347514 8195 353714 122064
rect 354494 8195 354734 122064
rect 355514 8195 361714 122064
rect 362494 121984 369714 122064
rect 370494 121984 378734 122064
rect 362494 8195 362734 121984
rect 363514 8195 369714 121984
rect 370494 8195 370734 121984
rect 371514 121940 378734 121984
rect 371514 8195 377714 121940
rect 378494 8195 378734 121940
rect 379514 121940 386734 122064
rect 379514 8195 385714 121940
rect 386494 8195 386734 121940
rect 387514 8195 393714 122064
rect 394494 8195 394734 122064
rect 395514 8195 401714 122064
rect 402494 121984 409714 122064
rect 402494 8195 402734 121984
rect 403514 8195 409714 121984
rect 410494 8195 410734 122064
rect 411514 8195 417714 122064
rect 418494 8195 418734 122064
rect 419514 8195 425714 294677
rect 426494 8195 426734 294677
rect 427514 8195 433714 294677
rect 434494 8195 434734 294677
rect 435514 8195 437125 294677
<< metal5 >>
rect 1056 291886 438888 292506
rect 1056 290866 438888 291486
rect 1056 283886 438888 284506
rect 1056 282866 438888 283486
rect 1056 275886 438888 276506
rect 1056 274866 438888 275486
rect 1056 267886 438888 268506
rect 1056 266866 438888 267486
rect 1056 259886 438888 260506
rect 1056 258866 438888 259486
rect 1056 251886 438888 252506
rect 1056 250866 438888 251486
rect 1056 243886 438888 244506
rect 1056 242866 438888 243486
rect 1056 235886 438888 236506
rect 1056 234866 438888 235486
rect 1056 227886 438888 228506
rect 1056 226866 438888 227486
rect 1056 219886 438888 220506
rect 1056 218866 438888 219486
rect 1056 211886 438888 212506
rect 1056 210866 438888 211486
rect 1056 203886 438888 204506
rect 1056 202866 438888 203486
rect 1056 195886 438888 196506
rect 1056 194866 438888 195486
rect 1056 187886 438888 188506
rect 1056 186866 438888 187486
rect 1056 179886 438888 180506
rect 1056 178866 438888 179486
rect 1056 171886 438888 172506
rect 1056 170866 438888 171486
rect 1056 163886 438888 164506
rect 1056 162866 438888 163486
rect 1056 155886 438888 156506
rect 1056 154866 438888 155486
rect 1056 147886 438888 148506
rect 1056 146866 438888 147486
rect 1056 139886 438888 140506
rect 1056 138866 438888 139486
rect 1056 131886 438888 132506
rect 1056 130866 438888 131486
rect 1056 123886 438888 124506
rect 1056 122866 438888 123486
rect 1056 115886 438888 116506
rect 1056 114866 438888 115486
rect 1056 107886 438888 108506
rect 1056 106866 438888 107486
rect 1056 99886 438888 100506
rect 1056 98866 438888 99486
rect 1056 91886 438888 92506
rect 1056 90866 438888 91486
rect 1056 83886 438888 84506
rect 1056 82866 438888 83486
rect 1056 75886 438888 76506
rect 1056 74866 438888 75486
rect 1056 67886 438888 68506
rect 1056 66866 438888 67486
rect 1056 59886 438888 60506
rect 1056 58866 438888 59486
rect 1056 51886 438888 52506
rect 1056 50866 438888 51486
rect 1056 43886 438888 44506
rect 1056 42866 438888 43486
rect 1056 35886 438888 36506
rect 1056 34866 438888 35486
rect 1056 27886 438888 28506
rect 1056 26866 438888 27486
rect 1056 19886 438888 20506
rect 1056 18866 438888 19486
rect 1056 11886 438888 12506
rect 1056 10866 438888 11486
rect 1056 3886 438888 4506
rect 1056 2866 438888 3486
<< obsm5 >>
rect 17780 156826 418300 162340
rect 17780 148826 418300 154546
rect 17780 140826 418300 146546
rect 17780 132826 418300 138546
rect 17780 124826 418300 130546
rect 17780 116826 418300 122546
rect 17780 108826 418300 114546
rect 17780 100826 418300 106546
rect 17780 92826 418300 98546
rect 17780 84826 418300 90546
rect 17780 76826 418300 82546
rect 17780 68826 418300 74546
rect 17780 60826 418300 66546
rect 17780 52826 418300 58546
rect 17780 44826 418300 50546
rect 17780 41660 418300 42546
<< labels >>
rlabel metal4 s 2814 2128 3434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 10814 2128 11434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 18814 2128 19434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 18814 209324 19434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 26814 2128 27434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 26814 209324 27434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 34814 2128 35434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 34814 209324 35434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42814 2128 43434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42814 209324 43434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50814 2128 51434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50814 209448 51434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58814 2128 59434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58814 209324 59434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66814 2128 67434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66814 209324 67434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 74814 2128 75434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 74814 209324 75434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 82814 2128 83434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 82814 209324 83434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 90814 2128 91434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 90814 209448 91434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 98814 2128 99434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 98814 209324 99434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 106814 2128 107434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 106814 209324 107434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 114814 2128 115434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 114814 209324 115434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 122814 2128 123434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 122814 209448 123434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 130814 2128 131434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 130814 209324 131434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138814 2128 139434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138814 209324 139434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 146814 2128 147434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 146814 209324 147434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 154814 2128 155434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 154814 209324 155434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 162814 2128 163434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 170814 2128 171434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 178814 2128 179434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 186814 2128 187434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 194814 2128 195434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 202814 2128 203434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 210814 2128 211434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218814 2128 219434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 226814 2128 227434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 234814 2128 235434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 242814 2128 243434 47231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 242814 53073 243434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 250814 2128 251434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 258814 2128 259434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 266814 2128 267434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 274814 2128 275434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 282814 2128 283434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 282814 209324 283434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 290814 2128 291434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 290814 209324 291434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298814 2128 299434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298814 209324 299434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 306814 2128 307434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 306814 209324 307434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 314814 2128 315434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 314814 209324 315434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 322814 2128 323434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 322814 209448 323434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 330814 2128 331434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 330814 209448 331434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 338814 2128 339434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 338814 209324 339434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 346814 2128 347434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 346814 209324 347434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 354814 2128 355434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 354814 209324 355434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 362814 2128 363434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 362814 209448 363434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 370814 2128 371434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 370814 209448 371434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 378814 2128 379434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 378814 209324 379434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 386814 2128 387434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 386814 209324 387434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 394814 2128 395434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 394814 209324 395434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 402814 2128 403434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 402814 209324 403434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 410814 2128 411434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 410814 209448 411434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 418814 2128 419434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 426814 2128 427434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 434814 2128 435434 297616 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3886 438888 4506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 11886 438888 12506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 19886 438888 20506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 27886 438888 28506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 35886 438888 36506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 43886 438888 44506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 51886 438888 52506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 59886 438888 60506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67886 438888 68506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 75886 438888 76506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 83886 438888 84506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 91886 438888 92506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 99886 438888 100506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 107886 438888 108506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 115886 438888 116506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 123886 438888 124506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 131886 438888 132506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 139886 438888 140506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 147886 438888 148506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 155886 438888 156506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 163886 438888 164506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 171886 438888 172506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 179886 438888 180506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 187886 438888 188506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 195886 438888 196506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 203886 438888 204506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 211886 438888 212506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 219886 438888 220506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 227886 438888 228506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 235886 438888 236506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 243886 438888 244506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 251886 438888 252506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 259886 438888 260506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 267886 438888 268506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 275886 438888 276506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 283886 438888 284506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 291886 438888 292506 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9794 2128 10414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 17794 2128 18414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 17794 209324 18414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 25794 2128 26414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 25794 209324 26414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 33794 2128 34414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 33794 209324 34414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 41794 2128 42414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 41794 209324 42414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 49794 2128 50414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 49794 209324 50414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 57794 2128 58414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 57794 209392 58414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65794 2128 66414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65794 209392 66414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 209324 74414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 81794 2128 82414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 81794 209324 82414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 89794 2128 90414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 89794 209324 90414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 97794 2128 98414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 97794 209324 98414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 105794 2128 106414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 105794 209392 106414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 113794 2128 114414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 113794 209324 114414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 121794 2128 122414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 121794 209324 122414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 129794 2128 130414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 129794 209324 130414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137794 2128 138414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137794 209392 138414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 145794 2128 146414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 145794 209324 146414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 153794 2128 154414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 153794 209324 154414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 161794 2128 162414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 169794 2128 170414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 177794 2128 178414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 185794 2128 186414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 193794 2128 194414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 201794 2128 202414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 209794 2128 210414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217794 2128 218414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 225794 2128 226414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 233794 2128 234414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 241794 2128 242414 37900 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 241794 54788 242414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 249794 2128 250414 37900 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 249794 54788 250414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 257794 2128 258414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 265794 2128 266414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 273794 2128 274414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 281794 2128 282414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 281794 209324 282414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 289794 2128 290414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 289794 209324 290414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297794 2128 298414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297794 209324 298414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 305794 2128 306414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 305794 209324 306414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 313794 2128 314414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 313794 209324 314414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 321794 2128 322414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 321794 209324 322414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 329794 2128 330414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 329794 209324 330414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 337794 2128 338414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 337794 209392 338414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 345794 2128 346414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 345794 209392 346414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 353794 2128 354414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 353794 209324 354414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 361794 2128 362414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 361794 209324 362414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 369794 2128 370414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 369794 209324 370414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 377794 2128 378414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 377794 209392 378414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 385794 2128 386414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 385794 209392 386414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 393794 2128 394414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 393794 209324 394414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 401794 2128 402414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 401794 209324 402414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 409794 2128 410414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 409794 209324 410414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 417794 2128 418414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 417794 209324 418414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 425794 2128 426414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 433794 2128 434414 297616 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2866 438888 3486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 10866 438888 11486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 18866 438888 19486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 26866 438888 27486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 34866 438888 35486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 42866 438888 43486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 50866 438888 51486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 58866 438888 59486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66866 438888 67486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 74866 438888 75486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 82866 438888 83486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 90866 438888 91486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 98866 438888 99486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 106866 438888 107486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 114866 438888 115486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 122866 438888 123486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 130866 438888 131486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 138866 438888 139486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 146866 438888 147486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 154866 438888 155486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 162866 438888 163486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 170866 438888 171486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 178866 438888 179486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 186866 438888 187486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 194866 438888 195486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 202866 438888 203486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 210866 438888 211486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 218866 438888 219486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 226866 438888 227486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 234866 438888 235486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 242866 438888 243486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 250866 438888 251486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 258866 438888 259486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 266866 438888 267486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 274866 438888 275486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 282866 438888 283486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 290866 438888 291486 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 439520 8712 440000 8832 6 gpio_dm0[0]
port 3 nsew signal output
rlabel metal3 s 439520 204552 440000 204672 6 gpio_dm0[10]
port 4 nsew signal output
rlabel metal3 s 439520 224136 440000 224256 6 gpio_dm0[11]
port 5 nsew signal output
rlabel metal3 s 439520 243720 440000 243840 6 gpio_dm0[12]
port 6 nsew signal output
rlabel metal3 s 439520 263304 440000 263424 6 gpio_dm0[13]
port 7 nsew signal output
rlabel metal3 s 439520 282888 440000 283008 6 gpio_dm0[14]
port 8 nsew signal output
rlabel metal2 s 424322 299520 424378 300000 6 gpio_dm0[15]
port 9 nsew signal output
rlabel metal2 s 375746 299520 375802 300000 6 gpio_dm0[16]
port 10 nsew signal output
rlabel metal2 s 327170 299520 327226 300000 6 gpio_dm0[17]
port 11 nsew signal output
rlabel metal2 s 278594 299520 278650 300000 6 gpio_dm0[18]
port 12 nsew signal output
rlabel metal2 s 230018 299520 230074 300000 6 gpio_dm0[19]
port 13 nsew signal output
rlabel metal3 s 439520 28296 440000 28416 6 gpio_dm0[1]
port 14 nsew signal output
rlabel metal2 s 181442 299520 181498 300000 6 gpio_dm0[20]
port 15 nsew signal output
rlabel metal2 s 132866 299520 132922 300000 6 gpio_dm0[21]
port 16 nsew signal output
rlabel metal2 s 84290 299520 84346 300000 6 gpio_dm0[22]
port 17 nsew signal output
rlabel metal2 s 35714 299520 35770 300000 6 gpio_dm0[23]
port 18 nsew signal output
rlabel metal3 s 0 282888 480 283008 6 gpio_dm0[24]
port 19 nsew signal output
rlabel metal3 s 0 263304 480 263424 6 gpio_dm0[25]
port 20 nsew signal output
rlabel metal3 s 0 243720 480 243840 6 gpio_dm0[26]
port 21 nsew signal output
rlabel metal3 s 0 224136 480 224256 6 gpio_dm0[27]
port 22 nsew signal output
rlabel metal3 s 0 204552 480 204672 6 gpio_dm0[28]
port 23 nsew signal output
rlabel metal3 s 0 184968 480 185088 6 gpio_dm0[29]
port 24 nsew signal output
rlabel metal3 s 439520 47880 440000 48000 6 gpio_dm0[2]
port 25 nsew signal output
rlabel metal3 s 0 165384 480 165504 6 gpio_dm0[30]
port 26 nsew signal output
rlabel metal3 s 0 145800 480 145920 6 gpio_dm0[31]
port 27 nsew signal output
rlabel metal3 s 0 126216 480 126336 6 gpio_dm0[32]
port 28 nsew signal output
rlabel metal3 s 0 106632 480 106752 6 gpio_dm0[33]
port 29 nsew signal output
rlabel metal3 s 0 87048 480 87168 6 gpio_dm0[34]
port 30 nsew signal output
rlabel metal3 s 0 67464 480 67584 6 gpio_dm0[35]
port 31 nsew signal output
rlabel metal3 s 0 47880 480 48000 6 gpio_dm0[36]
port 32 nsew signal output
rlabel metal3 s 0 28296 480 28416 6 gpio_dm0[37]
port 33 nsew signal output
rlabel metal2 s 21178 0 21234 480 6 gpio_dm0[38]
port 34 nsew signal output
rlabel metal2 s 70858 0 70914 480 6 gpio_dm0[39]
port 35 nsew signal output
rlabel metal3 s 439520 67464 440000 67584 6 gpio_dm0[3]
port 36 nsew signal output
rlabel metal2 s 120538 0 120594 480 6 gpio_dm0[40]
port 37 nsew signal output
rlabel metal2 s 170218 0 170274 480 6 gpio_dm0[41]
port 38 nsew signal output
rlabel metal2 s 219898 0 219954 480 6 gpio_dm0[42]
port 39 nsew signal output
rlabel metal2 s 269578 0 269634 480 6 gpio_dm0[43]
port 40 nsew signal output
rlabel metal3 s 439520 87048 440000 87168 6 gpio_dm0[4]
port 41 nsew signal output
rlabel metal3 s 439520 106632 440000 106752 6 gpio_dm0[5]
port 42 nsew signal output
rlabel metal3 s 439520 126216 440000 126336 6 gpio_dm0[6]
port 43 nsew signal output
rlabel metal3 s 439520 145800 440000 145920 6 gpio_dm0[7]
port 44 nsew signal output
rlabel metal3 s 439520 165384 440000 165504 6 gpio_dm0[8]
port 45 nsew signal output
rlabel metal3 s 439520 184968 440000 185088 6 gpio_dm0[9]
port 46 nsew signal output
rlabel metal3 s 439520 7080 440000 7200 6 gpio_dm1[0]
port 47 nsew signal output
rlabel metal3 s 439520 202920 440000 203040 6 gpio_dm1[10]
port 48 nsew signal output
rlabel metal3 s 439520 222504 440000 222624 6 gpio_dm1[11]
port 49 nsew signal output
rlabel metal3 s 439520 242088 440000 242208 6 gpio_dm1[12]
port 50 nsew signal output
rlabel metal3 s 439520 261672 440000 261792 6 gpio_dm1[13]
port 51 nsew signal output
rlabel metal3 s 439520 281256 440000 281376 6 gpio_dm1[14]
port 52 nsew signal output
rlabel metal2 s 428370 299520 428426 300000 6 gpio_dm1[15]
port 53 nsew signal output
rlabel metal2 s 379794 299520 379850 300000 6 gpio_dm1[16]
port 54 nsew signal output
rlabel metal2 s 331218 299520 331274 300000 6 gpio_dm1[17]
port 55 nsew signal output
rlabel metal2 s 282642 299520 282698 300000 6 gpio_dm1[18]
port 56 nsew signal output
rlabel metal2 s 234066 299520 234122 300000 6 gpio_dm1[19]
port 57 nsew signal output
rlabel metal3 s 439520 26664 440000 26784 6 gpio_dm1[1]
port 58 nsew signal output
rlabel metal2 s 185490 299520 185546 300000 6 gpio_dm1[20]
port 59 nsew signal output
rlabel metal2 s 136914 299520 136970 300000 6 gpio_dm1[21]
port 60 nsew signal output
rlabel metal2 s 88338 299520 88394 300000 6 gpio_dm1[22]
port 61 nsew signal output
rlabel metal2 s 39762 299520 39818 300000 6 gpio_dm1[23]
port 62 nsew signal output
rlabel metal3 s 0 284520 480 284640 6 gpio_dm1[24]
port 63 nsew signal output
rlabel metal3 s 0 264936 480 265056 6 gpio_dm1[25]
port 64 nsew signal output
rlabel metal3 s 0 245352 480 245472 6 gpio_dm1[26]
port 65 nsew signal output
rlabel metal3 s 0 225768 480 225888 6 gpio_dm1[27]
port 66 nsew signal output
rlabel metal3 s 0 206184 480 206304 6 gpio_dm1[28]
port 67 nsew signal output
rlabel metal3 s 0 186600 480 186720 6 gpio_dm1[29]
port 68 nsew signal output
rlabel metal3 s 439520 46248 440000 46368 6 gpio_dm1[2]
port 69 nsew signal output
rlabel metal3 s 0 167016 480 167136 6 gpio_dm1[30]
port 70 nsew signal output
rlabel metal3 s 0 147432 480 147552 6 gpio_dm1[31]
port 71 nsew signal output
rlabel metal3 s 0 127848 480 127968 6 gpio_dm1[32]
port 72 nsew signal output
rlabel metal3 s 0 108264 480 108384 6 gpio_dm1[33]
port 73 nsew signal output
rlabel metal3 s 0 88680 480 88800 6 gpio_dm1[34]
port 74 nsew signal output
rlabel metal3 s 0 69096 480 69216 6 gpio_dm1[35]
port 75 nsew signal output
rlabel metal3 s 0 49512 480 49632 6 gpio_dm1[36]
port 76 nsew signal output
rlabel metal3 s 0 29928 480 30048 6 gpio_dm1[37]
port 77 nsew signal output
rlabel metal2 s 17038 0 17094 480 6 gpio_dm1[38]
port 78 nsew signal output
rlabel metal2 s 66718 0 66774 480 6 gpio_dm1[39]
port 79 nsew signal output
rlabel metal3 s 439520 65832 440000 65952 6 gpio_dm1[3]
port 80 nsew signal output
rlabel metal2 s 116398 0 116454 480 6 gpio_dm1[40]
port 81 nsew signal output
rlabel metal2 s 166078 0 166134 480 6 gpio_dm1[41]
port 82 nsew signal output
rlabel metal2 s 215758 0 215814 480 6 gpio_dm1[42]
port 83 nsew signal output
rlabel metal2 s 265438 0 265494 480 6 gpio_dm1[43]
port 84 nsew signal output
rlabel metal3 s 439520 85416 440000 85536 6 gpio_dm1[4]
port 85 nsew signal output
rlabel metal3 s 439520 105000 440000 105120 6 gpio_dm1[5]
port 86 nsew signal output
rlabel metal3 s 439520 124584 440000 124704 6 gpio_dm1[6]
port 87 nsew signal output
rlabel metal3 s 439520 144168 440000 144288 6 gpio_dm1[7]
port 88 nsew signal output
rlabel metal3 s 439520 163752 440000 163872 6 gpio_dm1[8]
port 89 nsew signal output
rlabel metal3 s 439520 183336 440000 183456 6 gpio_dm1[9]
port 90 nsew signal output
rlabel metal3 s 439520 11976 440000 12096 6 gpio_dm2[0]
port 91 nsew signal output
rlabel metal3 s 439520 207816 440000 207936 6 gpio_dm2[10]
port 92 nsew signal output
rlabel metal3 s 439520 227400 440000 227520 6 gpio_dm2[11]
port 93 nsew signal output
rlabel metal3 s 439520 246984 440000 247104 6 gpio_dm2[12]
port 94 nsew signal output
rlabel metal3 s 439520 266568 440000 266688 6 gpio_dm2[13]
port 95 nsew signal output
rlabel metal3 s 439520 286152 440000 286272 6 gpio_dm2[14]
port 96 nsew signal output
rlabel metal2 s 416226 299520 416282 300000 6 gpio_dm2[15]
port 97 nsew signal output
rlabel metal2 s 367650 299520 367706 300000 6 gpio_dm2[16]
port 98 nsew signal output
rlabel metal2 s 319074 299520 319130 300000 6 gpio_dm2[17]
port 99 nsew signal output
rlabel metal2 s 270498 299520 270554 300000 6 gpio_dm2[18]
port 100 nsew signal output
rlabel metal2 s 221922 299520 221978 300000 6 gpio_dm2[19]
port 101 nsew signal output
rlabel metal3 s 439520 31560 440000 31680 6 gpio_dm2[1]
port 102 nsew signal output
rlabel metal2 s 173346 299520 173402 300000 6 gpio_dm2[20]
port 103 nsew signal output
rlabel metal2 s 124770 299520 124826 300000 6 gpio_dm2[21]
port 104 nsew signal output
rlabel metal2 s 76194 299520 76250 300000 6 gpio_dm2[22]
port 105 nsew signal output
rlabel metal2 s 27618 299520 27674 300000 6 gpio_dm2[23]
port 106 nsew signal output
rlabel metal3 s 0 279624 480 279744 6 gpio_dm2[24]
port 107 nsew signal output
rlabel metal3 s 0 260040 480 260160 6 gpio_dm2[25]
port 108 nsew signal output
rlabel metal3 s 0 240456 480 240576 6 gpio_dm2[26]
port 109 nsew signal output
rlabel metal3 s 0 220872 480 220992 6 gpio_dm2[27]
port 110 nsew signal output
rlabel metal3 s 0 201288 480 201408 6 gpio_dm2[28]
port 111 nsew signal output
rlabel metal3 s 0 181704 480 181824 6 gpio_dm2[29]
port 112 nsew signal output
rlabel metal3 s 439520 51144 440000 51264 6 gpio_dm2[2]
port 113 nsew signal output
rlabel metal3 s 0 162120 480 162240 6 gpio_dm2[30]
port 114 nsew signal output
rlabel metal3 s 0 142536 480 142656 6 gpio_dm2[31]
port 115 nsew signal output
rlabel metal3 s 0 122952 480 123072 6 gpio_dm2[32]
port 116 nsew signal output
rlabel metal3 s 0 103368 480 103488 6 gpio_dm2[33]
port 117 nsew signal output
rlabel metal3 s 0 83784 480 83904 6 gpio_dm2[34]
port 118 nsew signal output
rlabel metal3 s 0 64200 480 64320 6 gpio_dm2[35]
port 119 nsew signal output
rlabel metal3 s 0 44616 480 44736 6 gpio_dm2[36]
port 120 nsew signal output
rlabel metal3 s 0 25032 480 25152 6 gpio_dm2[37]
port 121 nsew signal output
rlabel metal2 s 29458 0 29514 480 6 gpio_dm2[38]
port 122 nsew signal output
rlabel metal2 s 79138 0 79194 480 6 gpio_dm2[39]
port 123 nsew signal output
rlabel metal3 s 439520 70728 440000 70848 6 gpio_dm2[3]
port 124 nsew signal output
rlabel metal2 s 128818 0 128874 480 6 gpio_dm2[40]
port 125 nsew signal output
rlabel metal2 s 178498 0 178554 480 6 gpio_dm2[41]
port 126 nsew signal output
rlabel metal2 s 228178 0 228234 480 6 gpio_dm2[42]
port 127 nsew signal output
rlabel metal2 s 277858 0 277914 480 6 gpio_dm2[43]
port 128 nsew signal output
rlabel metal3 s 439520 90312 440000 90432 6 gpio_dm2[4]
port 129 nsew signal output
rlabel metal3 s 439520 109896 440000 110016 6 gpio_dm2[5]
port 130 nsew signal output
rlabel metal3 s 439520 129480 440000 129600 6 gpio_dm2[6]
port 131 nsew signal output
rlabel metal3 s 439520 149064 440000 149184 6 gpio_dm2[7]
port 132 nsew signal output
rlabel metal3 s 439520 168648 440000 168768 6 gpio_dm2[8]
port 133 nsew signal output
rlabel metal3 s 439520 188232 440000 188352 6 gpio_dm2[9]
port 134 nsew signal output
rlabel metal3 s 439520 16872 440000 16992 6 gpio_ib_mode_sel[0]
port 135 nsew signal output
rlabel metal3 s 439520 212712 440000 212832 6 gpio_ib_mode_sel[10]
port 136 nsew signal output
rlabel metal3 s 439520 232296 440000 232416 6 gpio_ib_mode_sel[11]
port 137 nsew signal output
rlabel metal3 s 439520 251880 440000 252000 6 gpio_ib_mode_sel[12]
port 138 nsew signal output
rlabel metal3 s 439520 271464 440000 271584 6 gpio_ib_mode_sel[13]
port 139 nsew signal output
rlabel metal3 s 439520 291048 440000 291168 6 gpio_ib_mode_sel[14]
port 140 nsew signal output
rlabel metal2 s 404082 299520 404138 300000 6 gpio_ib_mode_sel[15]
port 141 nsew signal output
rlabel metal2 s 355506 299520 355562 300000 6 gpio_ib_mode_sel[16]
port 142 nsew signal output
rlabel metal2 s 306930 299520 306986 300000 6 gpio_ib_mode_sel[17]
port 143 nsew signal output
rlabel metal2 s 258354 299520 258410 300000 6 gpio_ib_mode_sel[18]
port 144 nsew signal output
rlabel metal2 s 209778 299520 209834 300000 6 gpio_ib_mode_sel[19]
port 145 nsew signal output
rlabel metal3 s 439520 36456 440000 36576 6 gpio_ib_mode_sel[1]
port 146 nsew signal output
rlabel metal2 s 161202 299520 161258 300000 6 gpio_ib_mode_sel[20]
port 147 nsew signal output
rlabel metal2 s 112626 299520 112682 300000 6 gpio_ib_mode_sel[21]
port 148 nsew signal output
rlabel metal2 s 64050 299520 64106 300000 6 gpio_ib_mode_sel[22]
port 149 nsew signal output
rlabel metal2 s 15474 299520 15530 300000 6 gpio_ib_mode_sel[23]
port 150 nsew signal output
rlabel metal3 s 0 274728 480 274848 6 gpio_ib_mode_sel[24]
port 151 nsew signal output
rlabel metal3 s 0 255144 480 255264 6 gpio_ib_mode_sel[25]
port 152 nsew signal output
rlabel metal3 s 0 235560 480 235680 6 gpio_ib_mode_sel[26]
port 153 nsew signal output
rlabel metal3 s 0 215976 480 216096 6 gpio_ib_mode_sel[27]
port 154 nsew signal output
rlabel metal3 s 0 196392 480 196512 6 gpio_ib_mode_sel[28]
port 155 nsew signal output
rlabel metal3 s 0 176808 480 176928 6 gpio_ib_mode_sel[29]
port 156 nsew signal output
rlabel metal3 s 439520 56040 440000 56160 6 gpio_ib_mode_sel[2]
port 157 nsew signal output
rlabel metal3 s 0 157224 480 157344 6 gpio_ib_mode_sel[30]
port 158 nsew signal output
rlabel metal3 s 0 137640 480 137760 6 gpio_ib_mode_sel[31]
port 159 nsew signal output
rlabel metal3 s 0 118056 480 118176 6 gpio_ib_mode_sel[32]
port 160 nsew signal output
rlabel metal3 s 0 98472 480 98592 6 gpio_ib_mode_sel[33]
port 161 nsew signal output
rlabel metal3 s 0 78888 480 79008 6 gpio_ib_mode_sel[34]
port 162 nsew signal output
rlabel metal3 s 0 59304 480 59424 6 gpio_ib_mode_sel[35]
port 163 nsew signal output
rlabel metal3 s 0 39720 480 39840 6 gpio_ib_mode_sel[36]
port 164 nsew signal output
rlabel metal3 s 0 20136 480 20256 6 gpio_ib_mode_sel[37]
port 165 nsew signal output
rlabel metal2 s 41878 0 41934 480 6 gpio_ib_mode_sel[38]
port 166 nsew signal output
rlabel metal2 s 91558 0 91614 480 6 gpio_ib_mode_sel[39]
port 167 nsew signal output
rlabel metal3 s 439520 75624 440000 75744 6 gpio_ib_mode_sel[3]
port 168 nsew signal output
rlabel metal2 s 141238 0 141294 480 6 gpio_ib_mode_sel[40]
port 169 nsew signal output
rlabel metal2 s 190918 0 190974 480 6 gpio_ib_mode_sel[41]
port 170 nsew signal output
rlabel metal2 s 240598 0 240654 480 6 gpio_ib_mode_sel[42]
port 171 nsew signal output
rlabel metal2 s 290278 0 290334 480 6 gpio_ib_mode_sel[43]
port 172 nsew signal output
rlabel metal3 s 439520 95208 440000 95328 6 gpio_ib_mode_sel[4]
port 173 nsew signal output
rlabel metal3 s 439520 114792 440000 114912 6 gpio_ib_mode_sel[5]
port 174 nsew signal output
rlabel metal3 s 439520 134376 440000 134496 6 gpio_ib_mode_sel[6]
port 175 nsew signal output
rlabel metal3 s 439520 153960 440000 154080 6 gpio_ib_mode_sel[7]
port 176 nsew signal output
rlabel metal3 s 439520 173544 440000 173664 6 gpio_ib_mode_sel[8]
port 177 nsew signal output
rlabel metal3 s 439520 193128 440000 193248 6 gpio_ib_mode_sel[9]
port 178 nsew signal output
rlabel metal3 s 439520 10344 440000 10464 6 gpio_ieb[0]
port 179 nsew signal output
rlabel metal3 s 439520 206184 440000 206304 6 gpio_ieb[10]
port 180 nsew signal output
rlabel metal3 s 439520 225768 440000 225888 6 gpio_ieb[11]
port 181 nsew signal output
rlabel metal3 s 439520 245352 440000 245472 6 gpio_ieb[12]
port 182 nsew signal output
rlabel metal3 s 439520 264936 440000 265056 6 gpio_ieb[13]
port 183 nsew signal output
rlabel metal3 s 439520 284520 440000 284640 6 gpio_ieb[14]
port 184 nsew signal output
rlabel metal2 s 420274 299520 420330 300000 6 gpio_ieb[15]
port 185 nsew signal output
rlabel metal2 s 371698 299520 371754 300000 6 gpio_ieb[16]
port 186 nsew signal output
rlabel metal2 s 323122 299520 323178 300000 6 gpio_ieb[17]
port 187 nsew signal output
rlabel metal2 s 274546 299520 274602 300000 6 gpio_ieb[18]
port 188 nsew signal output
rlabel metal2 s 225970 299520 226026 300000 6 gpio_ieb[19]
port 189 nsew signal output
rlabel metal3 s 439520 29928 440000 30048 6 gpio_ieb[1]
port 190 nsew signal output
rlabel metal2 s 177394 299520 177450 300000 6 gpio_ieb[20]
port 191 nsew signal output
rlabel metal2 s 128818 299520 128874 300000 6 gpio_ieb[21]
port 192 nsew signal output
rlabel metal2 s 80242 299520 80298 300000 6 gpio_ieb[22]
port 193 nsew signal output
rlabel metal2 s 31666 299520 31722 300000 6 gpio_ieb[23]
port 194 nsew signal output
rlabel metal3 s 0 281256 480 281376 6 gpio_ieb[24]
port 195 nsew signal output
rlabel metal3 s 0 261672 480 261792 6 gpio_ieb[25]
port 196 nsew signal output
rlabel metal3 s 0 242088 480 242208 6 gpio_ieb[26]
port 197 nsew signal output
rlabel metal3 s 0 222504 480 222624 6 gpio_ieb[27]
port 198 nsew signal output
rlabel metal3 s 0 202920 480 203040 6 gpio_ieb[28]
port 199 nsew signal output
rlabel metal3 s 0 183336 480 183456 6 gpio_ieb[29]
port 200 nsew signal output
rlabel metal3 s 439520 49512 440000 49632 6 gpio_ieb[2]
port 201 nsew signal output
rlabel metal3 s 0 163752 480 163872 6 gpio_ieb[30]
port 202 nsew signal output
rlabel metal3 s 0 144168 480 144288 6 gpio_ieb[31]
port 203 nsew signal output
rlabel metal3 s 0 124584 480 124704 6 gpio_ieb[32]
port 204 nsew signal output
rlabel metal3 s 0 105000 480 105120 6 gpio_ieb[33]
port 205 nsew signal output
rlabel metal3 s 0 85416 480 85536 6 gpio_ieb[34]
port 206 nsew signal output
rlabel metal3 s 0 65832 480 65952 6 gpio_ieb[35]
port 207 nsew signal output
rlabel metal3 s 0 46248 480 46368 6 gpio_ieb[36]
port 208 nsew signal output
rlabel metal3 s 0 26664 480 26784 6 gpio_ieb[37]
port 209 nsew signal output
rlabel metal2 s 25318 0 25374 480 6 gpio_ieb[38]
port 210 nsew signal output
rlabel metal2 s 74998 0 75054 480 6 gpio_ieb[39]
port 211 nsew signal output
rlabel metal3 s 439520 69096 440000 69216 6 gpio_ieb[3]
port 212 nsew signal output
rlabel metal2 s 124678 0 124734 480 6 gpio_ieb[40]
port 213 nsew signal output
rlabel metal2 s 174358 0 174414 480 6 gpio_ieb[41]
port 214 nsew signal output
rlabel metal2 s 224038 0 224094 480 6 gpio_ieb[42]
port 215 nsew signal output
rlabel metal2 s 273718 0 273774 480 6 gpio_ieb[43]
port 216 nsew signal output
rlabel metal3 s 439520 88680 440000 88800 6 gpio_ieb[4]
port 217 nsew signal output
rlabel metal3 s 439520 108264 440000 108384 6 gpio_ieb[5]
port 218 nsew signal output
rlabel metal3 s 439520 127848 440000 127968 6 gpio_ieb[6]
port 219 nsew signal output
rlabel metal3 s 439520 147432 440000 147552 6 gpio_ieb[7]
port 220 nsew signal output
rlabel metal3 s 439520 167016 440000 167136 6 gpio_ieb[8]
port 221 nsew signal output
rlabel metal3 s 439520 186600 440000 186720 6 gpio_ieb[9]
port 222 nsew signal output
rlabel metal3 s 439520 3816 440000 3936 6 gpio_in[0]
port 223 nsew signal input
rlabel metal3 s 439520 199656 440000 199776 6 gpio_in[10]
port 224 nsew signal input
rlabel metal3 s 439520 219240 440000 219360 6 gpio_in[11]
port 225 nsew signal input
rlabel metal3 s 439520 238824 440000 238944 6 gpio_in[12]
port 226 nsew signal input
rlabel metal3 s 439520 258408 440000 258528 6 gpio_in[13]
port 227 nsew signal input
rlabel metal3 s 439520 277992 440000 278112 6 gpio_in[14]
port 228 nsew signal input
rlabel metal2 s 436466 299520 436522 300000 6 gpio_in[15]
port 229 nsew signal input
rlabel metal2 s 387890 299520 387946 300000 6 gpio_in[16]
port 230 nsew signal input
rlabel metal2 s 339314 299520 339370 300000 6 gpio_in[17]
port 231 nsew signal input
rlabel metal2 s 290738 299520 290794 300000 6 gpio_in[18]
port 232 nsew signal input
rlabel metal2 s 242162 299520 242218 300000 6 gpio_in[19]
port 233 nsew signal input
rlabel metal3 s 439520 23400 440000 23520 6 gpio_in[1]
port 234 nsew signal input
rlabel metal2 s 193586 299520 193642 300000 6 gpio_in[20]
port 235 nsew signal input
rlabel metal2 s 145010 299520 145066 300000 6 gpio_in[21]
port 236 nsew signal input
rlabel metal2 s 96434 299520 96490 300000 6 gpio_in[22]
port 237 nsew signal input
rlabel metal2 s 47858 299520 47914 300000 6 gpio_in[23]
port 238 nsew signal input
rlabel metal3 s 0 287784 480 287904 6 gpio_in[24]
port 239 nsew signal input
rlabel metal3 s 0 268200 480 268320 6 gpio_in[25]
port 240 nsew signal input
rlabel metal3 s 0 248616 480 248736 6 gpio_in[26]
port 241 nsew signal input
rlabel metal3 s 0 229032 480 229152 6 gpio_in[27]
port 242 nsew signal input
rlabel metal3 s 0 209448 480 209568 6 gpio_in[28]
port 243 nsew signal input
rlabel metal3 s 0 189864 480 189984 6 gpio_in[29]
port 244 nsew signal input
rlabel metal3 s 439520 42984 440000 43104 6 gpio_in[2]
port 245 nsew signal input
rlabel metal3 s 0 170280 480 170400 6 gpio_in[30]
port 246 nsew signal input
rlabel metal3 s 0 150696 480 150816 6 gpio_in[31]
port 247 nsew signal input
rlabel metal3 s 0 131112 480 131232 6 gpio_in[32]
port 248 nsew signal input
rlabel metal3 s 0 111528 480 111648 6 gpio_in[33]
port 249 nsew signal input
rlabel metal3 s 0 91944 480 92064 6 gpio_in[34]
port 250 nsew signal input
rlabel metal3 s 0 72360 480 72480 6 gpio_in[35]
port 251 nsew signal input
rlabel metal3 s 0 52776 480 52896 6 gpio_in[36]
port 252 nsew signal input
rlabel metal3 s 0 33192 480 33312 6 gpio_in[37]
port 253 nsew signal input
rlabel metal2 s 8758 0 8814 480 6 gpio_in[38]
port 254 nsew signal input
rlabel metal2 s 58438 0 58494 480 6 gpio_in[39]
port 255 nsew signal input
rlabel metal3 s 439520 62568 440000 62688 6 gpio_in[3]
port 256 nsew signal input
rlabel metal2 s 108118 0 108174 480 6 gpio_in[40]
port 257 nsew signal input
rlabel metal2 s 157798 0 157854 480 6 gpio_in[41]
port 258 nsew signal input
rlabel metal2 s 207478 0 207534 480 6 gpio_in[42]
port 259 nsew signal input
rlabel metal2 s 257158 0 257214 480 6 gpio_in[43]
port 260 nsew signal input
rlabel metal3 s 439520 82152 440000 82272 6 gpio_in[4]
port 261 nsew signal input
rlabel metal3 s 439520 101736 440000 101856 6 gpio_in[5]
port 262 nsew signal input
rlabel metal3 s 439520 121320 440000 121440 6 gpio_in[6]
port 263 nsew signal input
rlabel metal3 s 439520 140904 440000 141024 6 gpio_in[7]
port 264 nsew signal input
rlabel metal3 s 439520 160488 440000 160608 6 gpio_in[8]
port 265 nsew signal input
rlabel metal3 s 439520 180072 440000 180192 6 gpio_in[9]
port 266 nsew signal input
rlabel metal3 s 439520 20136 440000 20256 6 gpio_loopback_one[0]
port 267 nsew signal input
rlabel metal3 s 439520 215976 440000 216096 6 gpio_loopback_one[10]
port 268 nsew signal input
rlabel metal3 s 439520 235560 440000 235680 6 gpio_loopback_one[11]
port 269 nsew signal input
rlabel metal3 s 439520 255144 440000 255264 6 gpio_loopback_one[12]
port 270 nsew signal input
rlabel metal3 s 439520 274728 440000 274848 6 gpio_loopback_one[13]
port 271 nsew signal input
rlabel metal3 s 439520 294312 440000 294432 6 gpio_loopback_one[14]
port 272 nsew signal input
rlabel metal2 s 395986 299520 396042 300000 6 gpio_loopback_one[15]
port 273 nsew signal input
rlabel metal2 s 347410 299520 347466 300000 6 gpio_loopback_one[16]
port 274 nsew signal input
rlabel metal2 s 298834 299520 298890 300000 6 gpio_loopback_one[17]
port 275 nsew signal input
rlabel metal2 s 250258 299520 250314 300000 6 gpio_loopback_one[18]
port 276 nsew signal input
rlabel metal2 s 201682 299520 201738 300000 6 gpio_loopback_one[19]
port 277 nsew signal input
rlabel metal3 s 439520 39720 440000 39840 6 gpio_loopback_one[1]
port 278 nsew signal input
rlabel metal2 s 153106 299520 153162 300000 6 gpio_loopback_one[20]
port 279 nsew signal input
rlabel metal2 s 104530 299520 104586 300000 6 gpio_loopback_one[21]
port 280 nsew signal input
rlabel metal2 s 55954 299520 56010 300000 6 gpio_loopback_one[22]
port 281 nsew signal input
rlabel metal2 s 7378 299520 7434 300000 6 gpio_loopback_one[23]
port 282 nsew signal input
rlabel metal3 s 0 271464 480 271584 6 gpio_loopback_one[24]
port 283 nsew signal input
rlabel metal3 s 0 251880 480 252000 6 gpio_loopback_one[25]
port 284 nsew signal input
rlabel metal3 s 0 232296 480 232416 6 gpio_loopback_one[26]
port 285 nsew signal input
rlabel metal3 s 0 212712 480 212832 6 gpio_loopback_one[27]
port 286 nsew signal input
rlabel metal3 s 0 193128 480 193248 6 gpio_loopback_one[28]
port 287 nsew signal input
rlabel metal3 s 0 173544 480 173664 6 gpio_loopback_one[29]
port 288 nsew signal input
rlabel metal3 s 439520 59304 440000 59424 6 gpio_loopback_one[2]
port 289 nsew signal input
rlabel metal3 s 0 153960 480 154080 6 gpio_loopback_one[30]
port 290 nsew signal input
rlabel metal3 s 0 134376 480 134496 6 gpio_loopback_one[31]
port 291 nsew signal input
rlabel metal3 s 0 114792 480 114912 6 gpio_loopback_one[32]
port 292 nsew signal input
rlabel metal3 s 0 95208 480 95328 6 gpio_loopback_one[33]
port 293 nsew signal input
rlabel metal3 s 0 75624 480 75744 6 gpio_loopback_one[34]
port 294 nsew signal input
rlabel metal3 s 0 56040 480 56160 6 gpio_loopback_one[35]
port 295 nsew signal input
rlabel metal3 s 0 36456 480 36576 6 gpio_loopback_one[36]
port 296 nsew signal input
rlabel metal3 s 0 16872 480 16992 6 gpio_loopback_one[37]
port 297 nsew signal input
rlabel metal2 s 50158 0 50214 480 6 gpio_loopback_one[38]
port 298 nsew signal input
rlabel metal2 s 99838 0 99894 480 6 gpio_loopback_one[39]
port 299 nsew signal input
rlabel metal3 s 439520 78888 440000 79008 6 gpio_loopback_one[3]
port 300 nsew signal input
rlabel metal2 s 149518 0 149574 480 6 gpio_loopback_one[40]
port 301 nsew signal input
rlabel metal2 s 199198 0 199254 480 6 gpio_loopback_one[41]
port 302 nsew signal input
rlabel metal2 s 248878 0 248934 480 6 gpio_loopback_one[42]
port 303 nsew signal input
rlabel metal2 s 298558 0 298614 480 6 gpio_loopback_one[43]
port 304 nsew signal input
rlabel metal3 s 439520 98472 440000 98592 6 gpio_loopback_one[4]
port 305 nsew signal input
rlabel metal3 s 439520 118056 440000 118176 6 gpio_loopback_one[5]
port 306 nsew signal input
rlabel metal3 s 439520 137640 440000 137760 6 gpio_loopback_one[6]
port 307 nsew signal input
rlabel metal3 s 439520 157224 440000 157344 6 gpio_loopback_one[7]
port 308 nsew signal input
rlabel metal3 s 439520 176808 440000 176928 6 gpio_loopback_one[8]
port 309 nsew signal input
rlabel metal3 s 439520 196392 440000 196512 6 gpio_loopback_one[9]
port 310 nsew signal input
rlabel metal3 s 439520 21768 440000 21888 6 gpio_loopback_zero[0]
port 311 nsew signal input
rlabel metal3 s 439520 217608 440000 217728 6 gpio_loopback_zero[10]
port 312 nsew signal input
rlabel metal3 s 439520 237192 440000 237312 6 gpio_loopback_zero[11]
port 313 nsew signal input
rlabel metal3 s 439520 256776 440000 256896 6 gpio_loopback_zero[12]
port 314 nsew signal input
rlabel metal3 s 439520 276360 440000 276480 6 gpio_loopback_zero[13]
port 315 nsew signal input
rlabel metal3 s 439520 295944 440000 296064 6 gpio_loopback_zero[14]
port 316 nsew signal input
rlabel metal2 s 391938 299520 391994 300000 6 gpio_loopback_zero[15]
port 317 nsew signal input
rlabel metal2 s 343362 299520 343418 300000 6 gpio_loopback_zero[16]
port 318 nsew signal input
rlabel metal2 s 294786 299520 294842 300000 6 gpio_loopback_zero[17]
port 319 nsew signal input
rlabel metal2 s 246210 299520 246266 300000 6 gpio_loopback_zero[18]
port 320 nsew signal input
rlabel metal2 s 197634 299520 197690 300000 6 gpio_loopback_zero[19]
port 321 nsew signal input
rlabel metal3 s 439520 41352 440000 41472 6 gpio_loopback_zero[1]
port 322 nsew signal input
rlabel metal2 s 149058 299520 149114 300000 6 gpio_loopback_zero[20]
port 323 nsew signal input
rlabel metal2 s 100482 299520 100538 300000 6 gpio_loopback_zero[21]
port 324 nsew signal input
rlabel metal2 s 51906 299520 51962 300000 6 gpio_loopback_zero[22]
port 325 nsew signal input
rlabel metal2 s 3330 299520 3386 300000 6 gpio_loopback_zero[23]
port 326 nsew signal input
rlabel metal3 s 0 269832 480 269952 6 gpio_loopback_zero[24]
port 327 nsew signal input
rlabel metal3 s 0 250248 480 250368 6 gpio_loopback_zero[25]
port 328 nsew signal input
rlabel metal3 s 0 230664 480 230784 6 gpio_loopback_zero[26]
port 329 nsew signal input
rlabel metal3 s 0 211080 480 211200 6 gpio_loopback_zero[27]
port 330 nsew signal input
rlabel metal3 s 0 191496 480 191616 6 gpio_loopback_zero[28]
port 331 nsew signal input
rlabel metal3 s 0 171912 480 172032 6 gpio_loopback_zero[29]
port 332 nsew signal input
rlabel metal3 s 439520 60936 440000 61056 6 gpio_loopback_zero[2]
port 333 nsew signal input
rlabel metal3 s 0 152328 480 152448 6 gpio_loopback_zero[30]
port 334 nsew signal input
rlabel metal3 s 0 132744 480 132864 6 gpio_loopback_zero[31]
port 335 nsew signal input
rlabel metal3 s 0 113160 480 113280 6 gpio_loopback_zero[32]
port 336 nsew signal input
rlabel metal3 s 0 93576 480 93696 6 gpio_loopback_zero[33]
port 337 nsew signal input
rlabel metal3 s 0 73992 480 74112 6 gpio_loopback_zero[34]
port 338 nsew signal input
rlabel metal3 s 0 54408 480 54528 6 gpio_loopback_zero[35]
port 339 nsew signal input
rlabel metal3 s 0 34824 480 34944 6 gpio_loopback_zero[36]
port 340 nsew signal input
rlabel metal3 s 0 15240 480 15360 6 gpio_loopback_zero[37]
port 341 nsew signal input
rlabel metal2 s 54298 0 54354 480 6 gpio_loopback_zero[38]
port 342 nsew signal input
rlabel metal2 s 103978 0 104034 480 6 gpio_loopback_zero[39]
port 343 nsew signal input
rlabel metal3 s 439520 80520 440000 80640 6 gpio_loopback_zero[3]
port 344 nsew signal input
rlabel metal2 s 153658 0 153714 480 6 gpio_loopback_zero[40]
port 345 nsew signal input
rlabel metal2 s 203338 0 203394 480 6 gpio_loopback_zero[41]
port 346 nsew signal input
rlabel metal2 s 253018 0 253074 480 6 gpio_loopback_zero[42]
port 347 nsew signal input
rlabel metal2 s 302698 0 302754 480 6 gpio_loopback_zero[43]
port 348 nsew signal input
rlabel metal3 s 439520 100104 440000 100224 6 gpio_loopback_zero[4]
port 349 nsew signal input
rlabel metal3 s 439520 119688 440000 119808 6 gpio_loopback_zero[5]
port 350 nsew signal input
rlabel metal3 s 439520 139272 440000 139392 6 gpio_loopback_zero[6]
port 351 nsew signal input
rlabel metal3 s 439520 158856 440000 158976 6 gpio_loopback_zero[7]
port 352 nsew signal input
rlabel metal3 s 439520 178440 440000 178560 6 gpio_loopback_zero[8]
port 353 nsew signal input
rlabel metal3 s 439520 198024 440000 198144 6 gpio_loopback_zero[9]
port 354 nsew signal input
rlabel metal3 s 439520 18504 440000 18624 6 gpio_oeb[0]
port 355 nsew signal output
rlabel metal3 s 439520 214344 440000 214464 6 gpio_oeb[10]
port 356 nsew signal output
rlabel metal3 s 439520 233928 440000 234048 6 gpio_oeb[11]
port 357 nsew signal output
rlabel metal3 s 439520 253512 440000 253632 6 gpio_oeb[12]
port 358 nsew signal output
rlabel metal3 s 439520 273096 440000 273216 6 gpio_oeb[13]
port 359 nsew signal output
rlabel metal3 s 439520 292680 440000 292800 6 gpio_oeb[14]
port 360 nsew signal output
rlabel metal2 s 400034 299520 400090 300000 6 gpio_oeb[15]
port 361 nsew signal output
rlabel metal2 s 351458 299520 351514 300000 6 gpio_oeb[16]
port 362 nsew signal output
rlabel metal2 s 302882 299520 302938 300000 6 gpio_oeb[17]
port 363 nsew signal output
rlabel metal2 s 254306 299520 254362 300000 6 gpio_oeb[18]
port 364 nsew signal output
rlabel metal2 s 205730 299520 205786 300000 6 gpio_oeb[19]
port 365 nsew signal output
rlabel metal3 s 439520 38088 440000 38208 6 gpio_oeb[1]
port 366 nsew signal output
rlabel metal2 s 157154 299520 157210 300000 6 gpio_oeb[20]
port 367 nsew signal output
rlabel metal2 s 108578 299520 108634 300000 6 gpio_oeb[21]
port 368 nsew signal output
rlabel metal2 s 60002 299520 60058 300000 6 gpio_oeb[22]
port 369 nsew signal output
rlabel metal2 s 11426 299520 11482 300000 6 gpio_oeb[23]
port 370 nsew signal output
rlabel metal3 s 0 273096 480 273216 6 gpio_oeb[24]
port 371 nsew signal output
rlabel metal3 s 0 253512 480 253632 6 gpio_oeb[25]
port 372 nsew signal output
rlabel metal3 s 0 233928 480 234048 6 gpio_oeb[26]
port 373 nsew signal output
rlabel metal3 s 0 214344 480 214464 6 gpio_oeb[27]
port 374 nsew signal output
rlabel metal3 s 0 194760 480 194880 6 gpio_oeb[28]
port 375 nsew signal output
rlabel metal3 s 0 175176 480 175296 6 gpio_oeb[29]
port 376 nsew signal output
rlabel metal3 s 439520 57672 440000 57792 6 gpio_oeb[2]
port 377 nsew signal output
rlabel metal3 s 0 155592 480 155712 6 gpio_oeb[30]
port 378 nsew signal output
rlabel metal3 s 0 136008 480 136128 6 gpio_oeb[31]
port 379 nsew signal output
rlabel metal3 s 0 116424 480 116544 6 gpio_oeb[32]
port 380 nsew signal output
rlabel metal3 s 0 96840 480 96960 6 gpio_oeb[33]
port 381 nsew signal output
rlabel metal3 s 0 77256 480 77376 6 gpio_oeb[34]
port 382 nsew signal output
rlabel metal3 s 0 57672 480 57792 6 gpio_oeb[35]
port 383 nsew signal output
rlabel metal3 s 0 38088 480 38208 6 gpio_oeb[36]
port 384 nsew signal output
rlabel metal3 s 0 18504 480 18624 6 gpio_oeb[37]
port 385 nsew signal output
rlabel metal2 s 46018 0 46074 480 6 gpio_oeb[38]
port 386 nsew signal output
rlabel metal2 s 95698 0 95754 480 6 gpio_oeb[39]
port 387 nsew signal output
rlabel metal3 s 439520 77256 440000 77376 6 gpio_oeb[3]
port 388 nsew signal output
rlabel metal2 s 145378 0 145434 480 6 gpio_oeb[40]
port 389 nsew signal output
rlabel metal2 s 195058 0 195114 480 6 gpio_oeb[41]
port 390 nsew signal output
rlabel metal2 s 244738 0 244794 480 6 gpio_oeb[42]
port 391 nsew signal output
rlabel metal2 s 294418 0 294474 480 6 gpio_oeb[43]
port 392 nsew signal output
rlabel metal3 s 439520 96840 440000 96960 6 gpio_oeb[4]
port 393 nsew signal output
rlabel metal3 s 439520 116424 440000 116544 6 gpio_oeb[5]
port 394 nsew signal output
rlabel metal3 s 439520 136008 440000 136128 6 gpio_oeb[6]
port 395 nsew signal output
rlabel metal3 s 439520 155592 440000 155712 6 gpio_oeb[7]
port 396 nsew signal output
rlabel metal3 s 439520 175176 440000 175296 6 gpio_oeb[8]
port 397 nsew signal output
rlabel metal3 s 439520 194760 440000 194880 6 gpio_oeb[9]
port 398 nsew signal output
rlabel metal3 s 439520 13608 440000 13728 6 gpio_out[0]
port 399 nsew signal output
rlabel metal3 s 439520 209448 440000 209568 6 gpio_out[10]
port 400 nsew signal output
rlabel metal3 s 439520 229032 440000 229152 6 gpio_out[11]
port 401 nsew signal output
rlabel metal3 s 439520 248616 440000 248736 6 gpio_out[12]
port 402 nsew signal output
rlabel metal3 s 439520 268200 440000 268320 6 gpio_out[13]
port 403 nsew signal output
rlabel metal3 s 439520 287784 440000 287904 6 gpio_out[14]
port 404 nsew signal output
rlabel metal2 s 412178 299520 412234 300000 6 gpio_out[15]
port 405 nsew signal output
rlabel metal2 s 363602 299520 363658 300000 6 gpio_out[16]
port 406 nsew signal output
rlabel metal2 s 315026 299520 315082 300000 6 gpio_out[17]
port 407 nsew signal output
rlabel metal2 s 266450 299520 266506 300000 6 gpio_out[18]
port 408 nsew signal output
rlabel metal2 s 217874 299520 217930 300000 6 gpio_out[19]
port 409 nsew signal output
rlabel metal3 s 439520 33192 440000 33312 6 gpio_out[1]
port 410 nsew signal output
rlabel metal2 s 169298 299520 169354 300000 6 gpio_out[20]
port 411 nsew signal output
rlabel metal2 s 120722 299520 120778 300000 6 gpio_out[21]
port 412 nsew signal output
rlabel metal2 s 72146 299520 72202 300000 6 gpio_out[22]
port 413 nsew signal output
rlabel metal2 s 23570 299520 23626 300000 6 gpio_out[23]
port 414 nsew signal output
rlabel metal3 s 0 277992 480 278112 6 gpio_out[24]
port 415 nsew signal output
rlabel metal3 s 0 258408 480 258528 6 gpio_out[25]
port 416 nsew signal output
rlabel metal3 s 0 238824 480 238944 6 gpio_out[26]
port 417 nsew signal output
rlabel metal3 s 0 219240 480 219360 6 gpio_out[27]
port 418 nsew signal output
rlabel metal3 s 0 199656 480 199776 6 gpio_out[28]
port 419 nsew signal output
rlabel metal3 s 0 180072 480 180192 6 gpio_out[29]
port 420 nsew signal output
rlabel metal3 s 439520 52776 440000 52896 6 gpio_out[2]
port 421 nsew signal output
rlabel metal3 s 0 160488 480 160608 6 gpio_out[30]
port 422 nsew signal output
rlabel metal3 s 0 140904 480 141024 6 gpio_out[31]
port 423 nsew signal output
rlabel metal3 s 0 121320 480 121440 6 gpio_out[32]
port 424 nsew signal output
rlabel metal3 s 0 101736 480 101856 6 gpio_out[33]
port 425 nsew signal output
rlabel metal3 s 0 82152 480 82272 6 gpio_out[34]
port 426 nsew signal output
rlabel metal3 s 0 62568 480 62688 6 gpio_out[35]
port 427 nsew signal output
rlabel metal3 s 0 42984 480 43104 6 gpio_out[36]
port 428 nsew signal output
rlabel metal3 s 0 23400 480 23520 6 gpio_out[37]
port 429 nsew signal output
rlabel metal2 s 33598 0 33654 480 6 gpio_out[38]
port 430 nsew signal output
rlabel metal2 s 83278 0 83334 480 6 gpio_out[39]
port 431 nsew signal output
rlabel metal3 s 439520 72360 440000 72480 6 gpio_out[3]
port 432 nsew signal output
rlabel metal2 s 132958 0 133014 480 6 gpio_out[40]
port 433 nsew signal output
rlabel metal2 s 182638 0 182694 480 6 gpio_out[41]
port 434 nsew signal output
rlabel metal2 s 232318 0 232374 480 6 gpio_out[42]
port 435 nsew signal output
rlabel metal2 s 281998 0 282054 480 6 gpio_out[43]
port 436 nsew signal output
rlabel metal3 s 439520 91944 440000 92064 6 gpio_out[4]
port 437 nsew signal output
rlabel metal3 s 439520 111528 440000 111648 6 gpio_out[5]
port 438 nsew signal output
rlabel metal3 s 439520 131112 440000 131232 6 gpio_out[6]
port 439 nsew signal output
rlabel metal3 s 439520 150696 440000 150816 6 gpio_out[7]
port 440 nsew signal output
rlabel metal3 s 439520 170280 440000 170400 6 gpio_out[8]
port 441 nsew signal output
rlabel metal3 s 439520 189864 440000 189984 6 gpio_out[9]
port 442 nsew signal output
rlabel metal3 s 439520 5448 440000 5568 6 gpio_slow_sel[0]
port 443 nsew signal output
rlabel metal3 s 439520 201288 440000 201408 6 gpio_slow_sel[10]
port 444 nsew signal output
rlabel metal3 s 439520 220872 440000 220992 6 gpio_slow_sel[11]
port 445 nsew signal output
rlabel metal3 s 439520 240456 440000 240576 6 gpio_slow_sel[12]
port 446 nsew signal output
rlabel metal3 s 439520 260040 440000 260160 6 gpio_slow_sel[13]
port 447 nsew signal output
rlabel metal3 s 439520 279624 440000 279744 6 gpio_slow_sel[14]
port 448 nsew signal output
rlabel metal2 s 432418 299520 432474 300000 6 gpio_slow_sel[15]
port 449 nsew signal output
rlabel metal2 s 383842 299520 383898 300000 6 gpio_slow_sel[16]
port 450 nsew signal output
rlabel metal2 s 335266 299520 335322 300000 6 gpio_slow_sel[17]
port 451 nsew signal output
rlabel metal2 s 286690 299520 286746 300000 6 gpio_slow_sel[18]
port 452 nsew signal output
rlabel metal2 s 238114 299520 238170 300000 6 gpio_slow_sel[19]
port 453 nsew signal output
rlabel metal3 s 439520 25032 440000 25152 6 gpio_slow_sel[1]
port 454 nsew signal output
rlabel metal2 s 189538 299520 189594 300000 6 gpio_slow_sel[20]
port 455 nsew signal output
rlabel metal2 s 140962 299520 141018 300000 6 gpio_slow_sel[21]
port 456 nsew signal output
rlabel metal2 s 92386 299520 92442 300000 6 gpio_slow_sel[22]
port 457 nsew signal output
rlabel metal2 s 43810 299520 43866 300000 6 gpio_slow_sel[23]
port 458 nsew signal output
rlabel metal3 s 0 286152 480 286272 6 gpio_slow_sel[24]
port 459 nsew signal output
rlabel metal3 s 0 266568 480 266688 6 gpio_slow_sel[25]
port 460 nsew signal output
rlabel metal3 s 0 246984 480 247104 6 gpio_slow_sel[26]
port 461 nsew signal output
rlabel metal3 s 0 227400 480 227520 6 gpio_slow_sel[27]
port 462 nsew signal output
rlabel metal3 s 0 207816 480 207936 6 gpio_slow_sel[28]
port 463 nsew signal output
rlabel metal3 s 0 188232 480 188352 6 gpio_slow_sel[29]
port 464 nsew signal output
rlabel metal3 s 439520 44616 440000 44736 6 gpio_slow_sel[2]
port 465 nsew signal output
rlabel metal3 s 0 168648 480 168768 6 gpio_slow_sel[30]
port 466 nsew signal output
rlabel metal3 s 0 149064 480 149184 6 gpio_slow_sel[31]
port 467 nsew signal output
rlabel metal3 s 0 129480 480 129600 6 gpio_slow_sel[32]
port 468 nsew signal output
rlabel metal3 s 0 109896 480 110016 6 gpio_slow_sel[33]
port 469 nsew signal output
rlabel metal3 s 0 90312 480 90432 6 gpio_slow_sel[34]
port 470 nsew signal output
rlabel metal3 s 0 70728 480 70848 6 gpio_slow_sel[35]
port 471 nsew signal output
rlabel metal3 s 0 51144 480 51264 6 gpio_slow_sel[36]
port 472 nsew signal output
rlabel metal3 s 0 31560 480 31680 6 gpio_slow_sel[37]
port 473 nsew signal output
rlabel metal2 s 12898 0 12954 480 6 gpio_slow_sel[38]
port 474 nsew signal output
rlabel metal2 s 62578 0 62634 480 6 gpio_slow_sel[39]
port 475 nsew signal output
rlabel metal3 s 439520 64200 440000 64320 6 gpio_slow_sel[3]
port 476 nsew signal output
rlabel metal2 s 112258 0 112314 480 6 gpio_slow_sel[40]
port 477 nsew signal output
rlabel metal2 s 161938 0 161994 480 6 gpio_slow_sel[41]
port 478 nsew signal output
rlabel metal2 s 211618 0 211674 480 6 gpio_slow_sel[42]
port 479 nsew signal output
rlabel metal2 s 261298 0 261354 480 6 gpio_slow_sel[43]
port 480 nsew signal output
rlabel metal3 s 439520 83784 440000 83904 6 gpio_slow_sel[4]
port 481 nsew signal output
rlabel metal3 s 439520 103368 440000 103488 6 gpio_slow_sel[5]
port 482 nsew signal output
rlabel metal3 s 439520 122952 440000 123072 6 gpio_slow_sel[6]
port 483 nsew signal output
rlabel metal3 s 439520 142536 440000 142656 6 gpio_slow_sel[7]
port 484 nsew signal output
rlabel metal3 s 439520 162120 440000 162240 6 gpio_slow_sel[8]
port 485 nsew signal output
rlabel metal3 s 439520 181704 440000 181824 6 gpio_slow_sel[9]
port 486 nsew signal output
rlabel metal3 s 439520 15240 440000 15360 6 gpio_vtrip_sel[0]
port 487 nsew signal output
rlabel metal3 s 439520 211080 440000 211200 6 gpio_vtrip_sel[10]
port 488 nsew signal output
rlabel metal3 s 439520 230664 440000 230784 6 gpio_vtrip_sel[11]
port 489 nsew signal output
rlabel metal3 s 439520 250248 440000 250368 6 gpio_vtrip_sel[12]
port 490 nsew signal output
rlabel metal3 s 439520 269832 440000 269952 6 gpio_vtrip_sel[13]
port 491 nsew signal output
rlabel metal3 s 439520 289416 440000 289536 6 gpio_vtrip_sel[14]
port 492 nsew signal output
rlabel metal2 s 408130 299520 408186 300000 6 gpio_vtrip_sel[15]
port 493 nsew signal output
rlabel metal2 s 359554 299520 359610 300000 6 gpio_vtrip_sel[16]
port 494 nsew signal output
rlabel metal2 s 310978 299520 311034 300000 6 gpio_vtrip_sel[17]
port 495 nsew signal output
rlabel metal2 s 262402 299520 262458 300000 6 gpio_vtrip_sel[18]
port 496 nsew signal output
rlabel metal2 s 213826 299520 213882 300000 6 gpio_vtrip_sel[19]
port 497 nsew signal output
rlabel metal3 s 439520 34824 440000 34944 6 gpio_vtrip_sel[1]
port 498 nsew signal output
rlabel metal2 s 165250 299520 165306 300000 6 gpio_vtrip_sel[20]
port 499 nsew signal output
rlabel metal2 s 116674 299520 116730 300000 6 gpio_vtrip_sel[21]
port 500 nsew signal output
rlabel metal2 s 68098 299520 68154 300000 6 gpio_vtrip_sel[22]
port 501 nsew signal output
rlabel metal2 s 19522 299520 19578 300000 6 gpio_vtrip_sel[23]
port 502 nsew signal output
rlabel metal3 s 0 276360 480 276480 6 gpio_vtrip_sel[24]
port 503 nsew signal output
rlabel metal3 s 0 256776 480 256896 6 gpio_vtrip_sel[25]
port 504 nsew signal output
rlabel metal3 s 0 237192 480 237312 6 gpio_vtrip_sel[26]
port 505 nsew signal output
rlabel metal3 s 0 217608 480 217728 6 gpio_vtrip_sel[27]
port 506 nsew signal output
rlabel metal3 s 0 198024 480 198144 6 gpio_vtrip_sel[28]
port 507 nsew signal output
rlabel metal3 s 0 178440 480 178560 6 gpio_vtrip_sel[29]
port 508 nsew signal output
rlabel metal3 s 439520 54408 440000 54528 6 gpio_vtrip_sel[2]
port 509 nsew signal output
rlabel metal3 s 0 158856 480 158976 6 gpio_vtrip_sel[30]
port 510 nsew signal output
rlabel metal3 s 0 139272 480 139392 6 gpio_vtrip_sel[31]
port 511 nsew signal output
rlabel metal3 s 0 119688 480 119808 6 gpio_vtrip_sel[32]
port 512 nsew signal output
rlabel metal3 s 0 100104 480 100224 6 gpio_vtrip_sel[33]
port 513 nsew signal output
rlabel metal3 s 0 80520 480 80640 6 gpio_vtrip_sel[34]
port 514 nsew signal output
rlabel metal3 s 0 60936 480 61056 6 gpio_vtrip_sel[35]
port 515 nsew signal output
rlabel metal3 s 0 41352 480 41472 6 gpio_vtrip_sel[36]
port 516 nsew signal output
rlabel metal3 s 0 21768 480 21888 6 gpio_vtrip_sel[37]
port 517 nsew signal output
rlabel metal2 s 37738 0 37794 480 6 gpio_vtrip_sel[38]
port 518 nsew signal output
rlabel metal2 s 87418 0 87474 480 6 gpio_vtrip_sel[39]
port 519 nsew signal output
rlabel metal3 s 439520 73992 440000 74112 6 gpio_vtrip_sel[3]
port 520 nsew signal output
rlabel metal2 s 137098 0 137154 480 6 gpio_vtrip_sel[40]
port 521 nsew signal output
rlabel metal2 s 186778 0 186834 480 6 gpio_vtrip_sel[41]
port 522 nsew signal output
rlabel metal2 s 236458 0 236514 480 6 gpio_vtrip_sel[42]
port 523 nsew signal output
rlabel metal2 s 286138 0 286194 480 6 gpio_vtrip_sel[43]
port 524 nsew signal output
rlabel metal3 s 439520 93576 440000 93696 6 gpio_vtrip_sel[4]
port 525 nsew signal output
rlabel metal3 s 439520 113160 440000 113280 6 gpio_vtrip_sel[5]
port 526 nsew signal output
rlabel metal3 s 439520 132744 440000 132864 6 gpio_vtrip_sel[6]
port 527 nsew signal output
rlabel metal3 s 439520 152328 440000 152448 6 gpio_vtrip_sel[7]
port 528 nsew signal output
rlabel metal3 s 439520 171912 440000 172032 6 gpio_vtrip_sel[8]
port 529 nsew signal output
rlabel metal3 s 439520 191496 440000 191616 6 gpio_vtrip_sel[9]
port 530 nsew signal output
rlabel metal2 s 306838 0 306894 480 6 mask_rev[0]
port 531 nsew signal input
rlabel metal2 s 348238 0 348294 480 6 mask_rev[10]
port 532 nsew signal input
rlabel metal2 s 352378 0 352434 480 6 mask_rev[11]
port 533 nsew signal input
rlabel metal2 s 356518 0 356574 480 6 mask_rev[12]
port 534 nsew signal input
rlabel metal2 s 360658 0 360714 480 6 mask_rev[13]
port 535 nsew signal input
rlabel metal2 s 364798 0 364854 480 6 mask_rev[14]
port 536 nsew signal input
rlabel metal2 s 368938 0 368994 480 6 mask_rev[15]
port 537 nsew signal input
rlabel metal2 s 373078 0 373134 480 6 mask_rev[16]
port 538 nsew signal input
rlabel metal2 s 377218 0 377274 480 6 mask_rev[17]
port 539 nsew signal input
rlabel metal2 s 381358 0 381414 480 6 mask_rev[18]
port 540 nsew signal input
rlabel metal2 s 385498 0 385554 480 6 mask_rev[19]
port 541 nsew signal input
rlabel metal2 s 310978 0 311034 480 6 mask_rev[1]
port 542 nsew signal input
rlabel metal2 s 389638 0 389694 480 6 mask_rev[20]
port 543 nsew signal input
rlabel metal2 s 393778 0 393834 480 6 mask_rev[21]
port 544 nsew signal input
rlabel metal2 s 397918 0 397974 480 6 mask_rev[22]
port 545 nsew signal input
rlabel metal2 s 402058 0 402114 480 6 mask_rev[23]
port 546 nsew signal input
rlabel metal2 s 406198 0 406254 480 6 mask_rev[24]
port 547 nsew signal input
rlabel metal2 s 410338 0 410394 480 6 mask_rev[25]
port 548 nsew signal input
rlabel metal2 s 414478 0 414534 480 6 mask_rev[26]
port 549 nsew signal input
rlabel metal2 s 418618 0 418674 480 6 mask_rev[27]
port 550 nsew signal input
rlabel metal2 s 422758 0 422814 480 6 mask_rev[28]
port 551 nsew signal input
rlabel metal2 s 426898 0 426954 480 6 mask_rev[29]
port 552 nsew signal input
rlabel metal2 s 315118 0 315174 480 6 mask_rev[2]
port 553 nsew signal input
rlabel metal2 s 431038 0 431094 480 6 mask_rev[30]
port 554 nsew signal input
rlabel metal2 s 435178 0 435234 480 6 mask_rev[31]
port 555 nsew signal input
rlabel metal2 s 319258 0 319314 480 6 mask_rev[3]
port 556 nsew signal input
rlabel metal2 s 323398 0 323454 480 6 mask_rev[4]
port 557 nsew signal input
rlabel metal2 s 327538 0 327594 480 6 mask_rev[5]
port 558 nsew signal input
rlabel metal2 s 331678 0 331734 480 6 mask_rev[6]
port 559 nsew signal input
rlabel metal2 s 335818 0 335874 480 6 mask_rev[7]
port 560 nsew signal input
rlabel metal2 s 339958 0 340014 480 6 mask_rev[8]
port 561 nsew signal input
rlabel metal2 s 344098 0 344154 480 6 mask_rev[9]
port 562 nsew signal input
rlabel metal3 s 0 13608 480 13728 6 por
port 563 nsew signal input
rlabel metal3 s 0 11976 480 12096 6 porb
port 564 nsew signal input
rlabel metal2 s 4618 0 4674 480 6 resetb
port 565 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 440000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 197701788
string GDS_FILE /home/hosni/caravel_openframe_project/openlane/picosoc/runs/23_08_08_17_02/results/signoff/picosoc.magic.gds
string GDS_START 18081820
<< end >>

